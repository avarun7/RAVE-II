module directory (

);

endmodule