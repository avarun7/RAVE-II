module cache_bank (

);

endmodule