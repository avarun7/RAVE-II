module directory (
    input clk,
    input rst, 


    //MEM_DATA_Q

    //MEM_INSTR_Q

    //I$_DATA_Q
    
    //I$_INSTR_Q

    //D$_DATA_Q

    //I$_INSTR_Q
    
);

endmodule