module d_split #(
    parameter OOO_TAG_SIZE = 10
    ) (
    
);
    
endmodule