module l2cache_TOP();

endmodule