module ras #(parameter XLEN=32, parameter DEPTH=128)(
    input clk, rst, valid_in,
    input push,
    input pop,

    output reg[XLEN-1:0] result,
    output reg       valid_out
);

initial begin
    
end

always @(posedge clk ) begin
    
end

endmodule