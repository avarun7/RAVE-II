module d_split #(
    parameter OOO_TAG_SIZE = 19
    ) (
    
);
    
endmodule