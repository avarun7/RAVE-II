module rob_TOP();

endmodule