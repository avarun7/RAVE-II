module dram_top #(parameter CL_SIZE = 128) (
    input clk,
    input rst,

    // I/O FROM INPUT QUEUES
    
    //EVEN SIDE
    //MEM_DATA_Q_in
    input[31:0] addr_in_mem_data_q_even,
    input [CL_SIZE-1:0] data_in_mem_data_q_even,
    input [2:0] operation_in_mem_data_q_even,
    input is_flush_in_mem_data_q_even,
    input alloc_in_mem_data_q_even,
    input [1:0] src_in_mem_data_q_even,
    input [1:0] dest_in_mem_data_q_even,

    output full_out_mem_data_q_even,
    
    //MEM_INSTR_Q_in
    input[31:0] addr_in_mem_instr_q_even,
    input [2:0] operation_in_mem_instr_q_even,
    input is_flush_in_mem_instr_q_even,
    input alloc_in_mem_instr_q_even,
    input [1:0] src_in_mem_instr_q_even,
    input [1:0] dest_in_mem_instr_q_even,

    output full_out_mem_instr_q_even,
    
    //ODD SIDE
    //MEM_DATA_Q_in
    input[31:0] addr_in_mem_data_q_odd,
    input [CL_SIZE-1:0] data_in_mem_data_q_odd,
    input [2:0] operation_in_mem_data_q_odd,
    input is_flush_in_mem_data_q_odd,
    input alloc_in_mem_data_q_odd,
    input [1:0] src_in_mem_data_q_odd,
    input [1:0] dest_in_mem_data_q_odd,

    output full_out_mem_data_q_odd,
    
    //MEM_INSTR_Q_in
    input[31:0] addr_in_mem_instr_q_odd,
    input [2:0] operation_in_mem_instr_q_odd,
    input is_flush_in_mem_instr_q_odd,
    input alloc_in_mem_instr_q_odd,
    input [1:0] src_in_mem_instr_q_odd,
    input [1:0] dest_in_mem_instr_q_odd,

    output full_out_mem_instr_q_odd,

    // I/O to OUTPUT QUEUES

    //EVEN SIDE
    //MEM_DATA_Q_out
    output [31:0] addr_out_mem_data_q_even,
    output [CL_SIZE-1:0] data_out_mem_data_q_even,
    output [2:0] operation_out_mem_data_q_even,
    output is_flush_out_mem_data_q_even,
    output alloc_out_mem_data_q_even,
    output [1:0] src_out_mem_data_q_even,
    output [1:0] dest_out_mem_data_q_even,

    input full_in_mem_data_q_even,

    //ODD SIDE
    //MEM_DATA_Q_out
    output [31:0] addr_out_mem_data_q_odd,
    output  [CL_SIZE-1:0] data_out_mem_data_q_odd,
    output  [2:0] operation_out_mem_data_q_odd,
    output  is_flush_out_mem_data_q_odd,
    output  alloc_out_mem_data_q_odd,
    output  [1:0] src_out_mem_data_q_odd,
    output  [1:0] dest_out_mem_data_q_odd,

    input full_in_mem_data_q_odd
);

       //MEM_DATA_Q_in
wire [31:0] bank_addr_in_mem_data_q_even;
wire  [CL_SIZE-1:0] bank_data_in_mem_data_q_even;
wire  [2:0] bank_operation_in_mem_data_q_even;
wire  bank_is_flush_in_mem_data_q_even;
wire  bank_valid_in_mem_data_q_even;
wire  [1:0] bank_src_in_mem_data_q_even;
wire  [1:0] bank_dest_in_mem_data_q_even;

wire [1:0] dealloc_even, dealloc_odd;
    //MEM_INSTR_Q_in
wire [31:0] bank_addr_in_mem_instr_q_even;
wire  [2:0] bank_operation_in_mem_instr_q_even;
wire  bank_is_flush_in_mem_instr_q_even;
wire  bank_valid_in_mem_instr_q_even;
wire  [1:0] bank_src_in_mem_instr_q_even;
wire  [1:0] bank_dest_in_mem_instr_q_even;
wire [CL_SIZE -1 : 0] bank_data_in_even, bank_data_in_odd;

data_q #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_data_q_even(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_data_q_even),
    .data_in(data_in_mem_data_q_even),
    .operation_in(operation_in_mem_data_q_even),
    .is_flush(is_flush_in_mem_data_q_even),
    .alloc(alloc_in_mem_data_q_even),
    .src(src_in_mem_data_q_even),
    .dest(dest_in_mem_data_q_even),
    //From reciever
    .dealloc(dealloc_even[1]),

    //output sender
    .full(full_out_mem_data_q_even),

    //output reciever
    .addr_out(bank_addr_in_mem_data_q_even),
    .data_out(bank_data_in_mem_data_q_even),
    .operation_out(bank_operation_in_mem_data_q_even),
    .valid(bank_valid_in_mem_data_q_even),
    .src_out(bank_src_in_mem_data_q_even),
    .dest_out(bank_dest_in_mem_data_q_even),
    .is_flush_out(bank_is_flush_in_mem_data_q_even)
);

instr_q  #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_instr_q_even(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_instr_q_even),
    .operation_in(operation_in_mem_instr_q_even),
    .is_flush(is_flush_in_mem_instr_q_even),
    .alloc(alloc_in_mem_instr_q_even),
    .src(src_in_mem_instr_q_even),
    .dest(dest_in_mem_instr_q_even),

    //From reciever
    .dealloc(dealloc_even[0]),

    //output sender
    .full(full_out_mem_instr_q_even),

    //output reciever
    .addr_out(bank_addr_in_mem_instr_q_even),
    .operation_out(bank_operation_in_mem_instr_q_even),
    .valid(bank_valid_in_mem_instr_q_even),
    .src_out(bank_src_in_mem_instr_q_even),
    .dest_out(bank_dest_in_mem_instr_q_even),
    .is_flush_out(bank_is_flush_in_mem_instr_q_even)
);
wire [31:0] bank_addr_in_even;
wire [2:0] bank_operation_in_even;
wire bank_valid_in_even;
// wire [CL_SIZE - 1:0] bank_data_in_even;
wire [1:0] bank_src_in_even;
wire [1:0] bank_dest_in_even;
wire bank_is_flush_in_even;

wire [31:0] bank_addr_in_odd;
wire [2:0] bank_operation_in_odd;
wire bank_valid_in_odd;
// wire [CL_SIZE - 1:0] bank_data_in_odd;
wire [1:0] bank_src_in_odd;
wire [1:0] bank_dest_in_odd;
wire bank_is_flush_in_odd;
queue_arbitrator #(.CL_SIZE(CL_SIZE), .Q_WIDTH(2)) queue_arb_even(
    .addr_in({
        bank_addr_in_mem_data_q_even,
        bank_addr_in_mem_instr_q_even
    }),
    .data_in({
        bank_data_in_mem_data_q_even,
        128'd0
    }),
    .operation_in({
        bank_operation_in_mem_data_q_even,
        bank_operation_in_mem_instr_q_even
    }), 
    .valid_in({
        bank_valid_in_mem_data_q_even,
        bank_valid_in_mem_instr_q_even
    }),
    .src_in({
        bank_src_in_mem_data_q_even,
        bank_src_in_mem_instr_q_even
    }),
    .dest_in({
        bank_dest_in_mem_data_q_even,
        bank_dest_in_mem_instr_q_even
    }),
    .is_flush_in({
        bank_is_flush_in_mem_data_q_even,
        bank_is_flush_in_mem_instr_q_even
    }),
    .stall_in(bank_stall_even),


    .addr_out(      bank_addr_in_even),
    .operation_out( bank_operation_in_even), 
    .valid_out(     bank_valid_in_even),
    .data_out(      bank_data_in_even),
    .src_out(       bank_src_in_even),
    .dest_out(      bank_dest_in_even),
    .is_flush_out(  bank_is_flush_in_even),

    .dealloc(dealloc_even)
);

dram_bank #(.CL_SIZE(CL_SIZE), .file_name(1)) db_even(
.rst(rst),
.clk(clk),

.addr_in(bank_addr_in_even),
.operation_in(bank_operation_in_even),
.valid_in(bank_valid_in_even),
.src_in(bank_src_in_even),
.dest_in(bank_dest_in_even),
.is_flush_in(bank_is_flush_in_even),
.data_in(bank_data_in_even),

.addr_out(addr_out_mem_data_q_even),
.operation_out(operation_out_mem_data_q_even),
.valid_out(alloc_out_mem_data_q_even),
.src_out(src_out_mem_data_q_even),
.dest_out(dest_out_mem_data_q_even),
.is_flush_out(is_flush_out_mem_data_q_even),
.data_out(data_out_mem_data_q_even),

.stall_out(bank_stall_even)
);
      //MEM_DATA_Q_in
wire [31:0] bank_addr_in_mem_data_q_odd;
wire  [CL_SIZE-1:0] bank_data_in_mem_data_q_odd;
wire  [2:0] bank_operation_in_mem_data_q_odd;
wire  bank_is_flush_in_mem_data_q_odd;
wire  bank_valid_in_mem_data_q_odd;
wire  [1:0] bank_src_in_mem_data_q_odd;
wire  [1:0] bank_dest_in_mem_data_q_odd;

    //MEM_INSTR_Q_in
wire [31:0] bank_addr_in_mem_instr_q_odd;
wire  [2:0] bank_operation_in_mem_instr_q_odd;
wire  bank_is_flush_in_mem_instr_q_odd;
wire  bank_valid_in_mem_instr_q_odd;
wire  [1:0] bank_src_in_mem_instr_q_odd;
wire  [1:0] bank_dest_in_mem_instr_q_odd;

data_q #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_data_q_odd(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_data_q_odd),
    .data_in(data_in_mem_data_q_odd),
    .operation_in(operation_in_mem_data_q_odd),
    .is_flush(is_flush_in_mem_data_q_odd),
    .alloc(alloc_in_mem_data_q_odd),
    .src(src_in_mem_data_q_odd),
    .dest(dest_in_mem_data_q_odd),
    //From reciever
    .dealloc(dealloc_odd[1]),

    //output sender
    .full(full_out_mem_data_q_odd),

    //output reciever
    .addr_out(bank_addr_in_mem_data_q_odd),
    .data_out(bank_data_in_mem_data_q_odd),
    .operation_out(bank_operation_in_mem_data_q_odd),
    .valid(bank_valid_in_mem_data_q_odd),
    .src_out(bank_src_in_mem_data_q_odd),
    .dest_out(bank_dest_in_mem_data_q_odd),
    .is_flush_out(bank_is_flush_in_mem_data_q_odd)
);

instr_q  #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_instr_q_odd(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_instr_q_odd),
    .operation_in(operation_in_mem_instr_q_odd),
    .is_flush(is_flush_in_mem_instr_q_odd),
    .alloc(alloc_in_mem_instr_q_odd),
    .src(src_in_mem_instr_q_odd),
    .dest(dest_in_mem_instr_q_odd),

    //From reciever
    .dealloc(dealloc_odd[0]),

    //output sender
    .full(full_out_mem_instr_q_odd),

    //output reciever
    .addr_out(bank_addr_in_mem_instr_q_odd),
    .operation_out(bank_operation_in_mem_instr_q_odd),
    .valid(bank_valid_in_mem_instr_q_odd),
    .src_out(bank_src_in_mem_instr_q_odd),
    .dest_out(bank_dest_in_mem_instr_q_odd),
    .is_flush_out(bank_is_flush_in_mem_instr_q_odd)
);
queue_arbitrator #(.CL_SIZE(CL_SIZE), .Q_WIDTH(2)) queue_arb_odd(
    .addr_in({
        bank_addr_in_mem_data_q_odd,
        bank_addr_in_mem_instr_q_odd
    }),
    .data_in({
        bank_data_in_mem_data_q_odd,
        128'd0
    }),
    .operation_in({
        bank_operation_in_mem_data_q_odd,
        bank_operation_in_mem_instr_q_odd
    }), 
    .valid_in({
        bank_valid_in_mem_data_q_odd,
        bank_valid_in_mem_instr_q_odd
    }),
    .src_in({
        bank_src_in_mem_data_q_odd,
        bank_src_in_mem_instr_q_odd
    }),
    .dest_in({
        bank_dest_in_mem_data_q_odd,
        bank_dest_in_mem_instr_q_odd
    }),
    .is_flush_in({
        bank_is_flush_in_mem_data_q_odd,
        bank_is_flush_in_mem_instr_q_odd
    }),

    .stall_in(bank_stall_odd),

    .addr_out(bank_addr_in_odd),
    .operation_out(bank_operation_in_odd), 
    .valid_out(bank_valid_in_odd),
    .data_out(bank_data_in_odd),
    .src_out(bank_src_in_odd),
    .dest_out(bank_dest_in_odd),
    .is_flush_out(bank_is_flush_in_odd),

    .dealloc(dealloc_odd)
);

dram_bank #(.CL_SIZE(128), .file_name(2)) db_odd(
.rst(rst),
.clk(clk),

.addr_in(bank_addr_in_odd),
.operation_in(bank_operation_in_odd),
.valid_in(bank_valid_in_odd),
.src_in(bank_src_in_odd),
.dest_in(bank_dest_in_odd),
.is_flush_in(bank_is_flush_in_odd),
.data_in(bank_data_in_odd),

.addr_out(addr_out_mem_data_q_odd),
.operation_out(operation_out_mem_data_q_odd),
.valid_out(alloc_out_mem_data_q_odd),
.src_out(src_out_mem_data_q_odd),
.dest_out(dest_out_mem_data_q_odd),
.is_flush_out(is_flush_out_mem_data_q_odd),
.data_out(data_out_mem_data_q_odd),

.stall_out(bank_stall_odd)
);


integer file;
  integer count = 0;
initial begin
    file = $fopen("MEM_FINAL.csv", "w");
    if (file == 0) begin
      $display("Error: Unable to open file.");
      $stop;
    end
    $fdisplay(file, "Little Endian - Smallest address on the right, largest address left\n");

    #100000
    $fdisplay(file, "0x0,0x%h_0x%h\n0x20,0x%h_0x%h\n0x40,0x%h_0x%h\n0x60,0x%h_0x%h\n0x80,0x%h_0x%h\n0xA0,0x%h_0x%h\n0xC0,0x%h_0x%h\n0xE0,0x%h_0x%h\n0x100,0x%h_0x%h\n0x120,0x%h_0x%h\n0x140,0x%h_0x%h\n0x160,0x%h_0x%h\n0x180,0x%h_0x%h\n0x1A0,0x%h_0x%h\n0x1C0,0x%h_0x%h\n0x1E0,0x%h_0x%h\n0x200,0x%h_0x%h\n0x220,0x%h_0x%h\n0x240,0x%h_0x%h\n0x260,0x%h_0x%h\n0x280,0x%h_0x%h\n0x2A0,0x%h_0x%h\n0x2C0,0x%h_0x%h\n0x2E0,0x%h_0x%h\n0x300,0x%h_0x%h\n0x320,0x%h_0x%h\n0x340,0x%h_0x%h\n0x360,0x%h_0x%h\n0x380,0x%h_0x%h\n0x3A0,0x%h_0x%h\n0x3C0,0x%h_0x%h\n0x3E0,0x%h_0x%h\n0x400,0x%h_0x%h\n0x420,0x%h_0x%h\n0x440,0x%h_0x%h\n0x460,0x%h_0x%h\n0x480,0x%h_0x%h\n0x4A0,0x%h_0x%h\n0x4C0,0x%h_0x%h\n0x4E0,0x%h_0x%h\n0x500,0x%h_0x%h\n0x520,0x%h_0x%h\n0x540,0x%h_0x%h\n0x560,0x%h_0x%h\n0x580,0x%h_0x%h\n0x5A0,0x%h_0x%h\n0x5C0,0x%h_0x%h\n0x5E0,0x%h_0x%h\n0x600,0x%h_0x%h\n0x620,0x%h_0x%h\n0x640,0x%h_0x%h\n0x660,0x%h_0x%h\n0x680,0x%h_0x%h\n0x6A0,0x%h_0x%h\n0x6C0,0x%h_0x%h\n0x6E0,0x%h_0x%h\n0x700,0x%h_0x%h\n0x720,0x%h_0x%h\n0x740,0x%h_0x%h\n0x760,0x%h_0x%h\n0x780,0x%h_0x%h\n0x7A0,0x%h_0x%h\n0x7C0,0x%h_0x%h\n0x7E0,0x%h_0x%h\n0x800,0x%h_0x%h\n0x820,0x%h_0x%h\n0x840,0x%h_0x%h\n0x860,0x%h_0x%h\n0x880,0x%h_0x%h\n0x8A0,0x%h_0x%h\n0x8C0,0x%h_0x%h\n0x8E0,0x%h_0x%h\n0x900,0x%h_0x%h\n0x920,0x%h_0x%h\n0x940,0x%h_0x%h\n0x960,0x%h_0x%h\n0x980,0x%h_0x%h\n0x9A0,0x%h_0x%h\n0x9C0,0x%h_0x%h\n0x9E0,0x%h_0x%h\n0xA00,0x%h_0x%h\n0xA20,0x%h_0x%h\n0xA40,0x%h_0x%h\n0xA60,0x%h_0x%h\n0xA80,0x%h_0x%h\n0xAA0,0x%h_0x%h\n0xAC0,0x%h_0x%h\n0xAE0,0x%h_0x%h\n0xB00,0x%h_0x%h\n0xB20,0x%h_0x%h\n0xB40,0x%h_0x%h\n0xB60,0x%h_0x%h\n0xB80,0x%h_0x%h\n0xBA0,0x%h_0x%h\n0xBC0,0x%h_0x%h\n0xBE0,0x%h_0x%h\n0xC00,0x%h_0x%h\n0xC20,0x%h_0x%h\n0xC40,0x%h_0x%h\n0xC60,0x%h_0x%h\n0xC80,0x%h_0x%h\n0xCA0,0x%h_0x%h\n0xCC0,0x%h_0x%h\n0xCE0,0x%h_0x%h\n0xD00,0x%h_0x%h\n0xD20,0x%h_0x%h\n0xD40,0x%h_0x%h\n0xD60,0x%h_0x%h\n0xD80,0x%h_0x%h\n0xDA0,0x%h_0x%h\n0xDC0,0x%h_0x%h\n0xDE0,0x%h_0x%h\n0xE00,0x%h_0x%h\n0xE20,0x%h_0x%h\n0xE40,0x%h_0x%h\n0xE60,0x%h_0x%h\n0xE80,0x%h_0x%h\n0xEA0,0x%h_0x%h\n0xEC0,0x%h_0x%h\n0xEE0,0x%h_0x%h\n0xF00,0x%h_0x%h\n0xF20,0x%h_0x%h\n0xF40,0x%h_0x%h\n0xF60,0x%h_0x%h\n0xF80,0x%h_0x%h\n0xFA0,0x%h_0x%h\n0xFC0,0x%h_0x%h\n0xFE0,0x%h_0x%h\n0x1000,0x%h_0x%h\n0x1020,0x%h_0x%h\n0x1040,0x%h_0x%h\n0x1060,0x%h_0x%h\n0x1080,0x%h_0x%h\n0x10A0,0x%h_0x%h\n0x10C0,0x%h_0x%h\n0x10E0,0x%h_0x%h\n0x1100,0x%h_0x%h\n0x1120,0x%h_0x%h\n0x1140,0x%h_0x%h\n0x1160,0x%h_0x%h\n0x1180,0x%h_0x%h\n0x11A0,0x%h_0x%h\n0x11C0,0x%h_0x%h\n0x11E0,0x%h_0x%h\n0x1200,0x%h_0x%h\n0x1220,0x%h_0x%h\n0x1240,0x%h_0x%h\n0x1260,0x%h_0x%h\n0x1280,0x%h_0x%h\n0x12A0,0x%h_0x%h\n0x12C0,0x%h_0x%h\n0x12E0,0x%h_0x%h\n0x1300,0x%h_0x%h\n0x1320,0x%h_0x%h\n0x1340,0x%h_0x%h\n0x1360,0x%h_0x%h\n0x1380,0x%h_0x%h\n0x13A0,0x%h_0x%h\n0x13C0,0x%h_0x%h\n0x13E0,0x%h_0x%h\n0x1400,0x%h_0x%h\n0x1420,0x%h_0x%h\n0x1440,0x%h_0x%h\n0x1460,0x%h_0x%h\n0x1480,0x%h_0x%h\n0x14A0,0x%h_0x%h\n0x14C0,0x%h_0x%h\n0x14E0,0x%h_0x%h\n0x1500,0x%h_0x%h\n0x1520,0x%h_0x%h\n0x1540,0x%h_0x%h\n0x1560,0x%h_0x%h\n0x1580,0x%h_0x%h\n0x15A0,0x%h_0x%h\n0x15C0,0x%h_0x%h\n0x15E0,0x%h_0x%h\n0x1600,0x%h_0x%h\n0x1620,0x%h_0x%h\n0x1640,0x%h_0x%h\n0x1660,0x%h_0x%h\n0x1680,0x%h_0x%h\n0x16A0,0x%h_0x%h\n0x16C0,0x%h_0x%h\n0x16E0,0x%h_0x%h\n0x1700,0x%h_0x%h\n0x1720,0x%h_0x%h\n0x1740,0x%h_0x%h\n0x1760,0x%h_0x%h\n0x1780,0x%h_0x%h\n0x17A0,0x%h_0x%h\n0x17C0,0x%h_0x%h\n0x17E0,0x%h_0x%h\n0x1800,0x%h_0x%h\n0x1820,0x%h_0x%h\n0x1840,0x%h_0x%h\n0x1860,0x%h_0x%h\n0x1880,0x%h_0x%h\n0x18A0,0x%h_0x%h\n0x18C0,0x%h_0x%h\n0x18E0,0x%h_0x%h\n0x1900,0x%h_0x%h\n0x1920,0x%h_0x%h\n0x1940,0x%h_0x%h\n0x1960,0x%h_0x%h\n0x1980,0x%h_0x%h\n0x19A0,0x%h_0x%h\n0x19C0,0x%h_0x%h\n0x19E0,0x%h_0x%h\n0x1A00,0x%h_0x%h\n0x1A20,0x%h_0x%h\n0x1A40,0x%h_0x%h\n0x1A60,0x%h_0x%h\n0x1A80,0x%h_0x%h\n0x1AA0,0x%h_0x%h\n0x1AC0,0x%h_0x%h\n0x1AE0,0x%h_0x%h\n0x1B00,0x%h_0x%h\n0x1B20,0x%h_0x%h\n0x1B40,0x%h_0x%h\n0x1B60,0x%h_0x%h\n0x1B80,0x%h_0x%h\n0x1BA0,0x%h_0x%h\n0x1BC0,0x%h_0x%h\n0x1BE0,0x%h_0x%h\n0x1C00,0x%h_0x%h\n0x1C20,0x%h_0x%h\n0x1C40,0x%h_0x%h\n0x1C60,0x%h_0x%h\n0x1C80,0x%h_0x%h\n0x1CA0,0x%h_0x%h\n0x1CC0,0x%h_0x%h\n0x1CE0,0x%h_0x%h\n0x1D00,0x%h_0x%h\n0x1D20,0x%h_0x%h\n0x1D40,0x%h_0x%h\n0x1D60,0x%h_0x%h\n0x1D80,0x%h_0x%h\n0x1DA0,0x%h_0x%h\n0x1DC0,0x%h_0x%h\n0x1DE0,0x%h_0x%h\n0x1E00,0x%h_0x%h\n0x1E20,0x%h_0x%h\n0x1E40,0x%h_0x%h\n0x1E60,0x%h_0x%h\n0x1E80,0x%h_0x%h\n0x1EA0,0x%h_0x%h\n0x1EC0,0x%h_0x%h\n0x1EE0,0x%h_0x%h\n0x1F00,0x%h_0x%h\n0x1F20,0x%h_0x%h\n0x1F40,0x%h_0x%h\n0x1F60,0x%h_0x%h\n0x1F80,0x%h_0x%h\n0x1FA0,0x%h_0x%h\n0x1FC0,0x%h_0x%h\n0x1FE0,0x%h_0x%h\n0x2000,0x%h_0x%h\n0x2020,0x%h_0x%h\n0x2040,0x%h_0x%h\n0x2060,0x%h_0x%h\n0x2080,0x%h_0x%h\n0x20A0,0x%h_0x%h\n0x20C0,0x%h_0x%h\n0x20E0,0x%h_0x%h\n0x2100,0x%h_0x%h\n0x2120,0x%h_0x%h\n0x2140,0x%h_0x%h\n0x2160,0x%h_0x%h\n0x2180,0x%h_0x%h\n0x21A0,0x%h_0x%h\n0x21C0,0x%h_0x%h\n0x21E0,0x%h_0x%h\n0x2200,0x%h_0x%h\n0x2220,0x%h_0x%h\n0x2240,0x%h_0x%h\n0x2260,0x%h_0x%h\n0x2280,0x%h_0x%h\n0x22A0,0x%h_0x%h\n0x22C0,0x%h_0x%h\n0x22E0,0x%h_0x%h\n0x2300,0x%h_0x%h\n0x2320,0x%h_0x%h\n0x2340,0x%h_0x%h\n0x2360,0x%h_0x%h\n0x2380,0x%h_0x%h\n0x23A0,0x%h_0x%h\n0x23C0,0x%h_0x%h\n0x23E0,0x%h_0x%h\n0x2400,0x%h_0x%h\n0x2420,0x%h_0x%h\n0x2440,0x%h_0x%h\n0x2460,0x%h_0x%h\n0x2480,0x%h_0x%h\n0x24A0,0x%h_0x%h\n0x24C0,0x%h_0x%h\n0x24E0,0x%h_0x%h\n0x2500,0x%h_0x%h\n0x2520,0x%h_0x%h\n0x2540,0x%h_0x%h\n0x2560,0x%h_0x%h\n0x2580,0x%h_0x%h\n0x25A0,0x%h_0x%h\n0x25C0,0x%h_0x%h\n0x25E0,0x%h_0x%h\n0x2600,0x%h_0x%h\n0x2620,0x%h_0x%h\n0x2640,0x%h_0x%h\n0x2660,0x%h_0x%h\n0x2680,0x%h_0x%h\n0x26A0,0x%h_0x%h\n0x26C0,0x%h_0x%h\n0x26E0,0x%h_0x%h\n0x2700,0x%h_0x%h\n0x2720,0x%h_0x%h\n0x2740,0x%h_0x%h\n0x2760,0x%h_0x%h\n0x2780,0x%h_0x%h\n0x27A0,0x%h_0x%h\n0x27C0,0x%h_0x%h\n0x27E0,0x%h_0x%h\n0x2800,0x%h_0x%h\n0x2820,0x%h_0x%h\n0x2840,0x%h_0x%h\n0x2860,0x%h_0x%h\n0x2880,0x%h_0x%h\n0x28A0,0x%h_0x%h\n0x28C0,0x%h_0x%h\n0x28E0,0x%h_0x%h\n0x2900,0x%h_0x%h\n0x2920,0x%h_0x%h\n0x2940,0x%h_0x%h\n0x2960,0x%h_0x%h\n0x2980,0x%h_0x%h\n0x29A0,0x%h_0x%h\n0x29C0,0x%h_0x%h\n0x29E0,0x%h_0x%h\n0x2A00,0x%h_0x%h\n0x2A20,0x%h_0x%h\n0x2A40,0x%h_0x%h\n0x2A60,0x%h_0x%h\n0x2A80,0x%h_0x%h\n0x2AA0,0x%h_0x%h\n0x2AC0,0x%h_0x%h\n0x2AE0,0x%h_0x%h\n0x2B00,0x%h_0x%h\n0x2B20,0x%h_0x%h\n0x2B40,0x%h_0x%h\n0x2B60,0x%h_0x%h\n0x2B80,0x%h_0x%h\n0x2BA0,0x%h_0x%h\n0x2BC0,0x%h_0x%h\n0x2BE0,0x%h_0x%h\n0x2C00,0x%h_0x%h\n0x2C20,0x%h_0x%h\n0x2C40,0x%h_0x%h\n0x2C60,0x%h_0x%h\n0x2C80,0x%h_0x%h\n0x2CA0,0x%h_0x%h\n0x2CC0,0x%h_0x%h\n0x2CE0,0x%h_0x%h\n0x2D00,0x%h_0x%h\n0x2D20,0x%h_0x%h\n0x2D40,0x%h_0x%h\n0x2D60,0x%h_0x%h\n0x2D80,0x%h_0x%h\n0x2DA0,0x%h_0x%h\n0x2DC0,0x%h_0x%h\n0x2DE0,0x%h_0x%h\n0x2E00,0x%h_0x%h\n0x2E20,0x%h_0x%h\n0x2E40,0x%h_0x%h\n0x2E60,0x%h_0x%h\n0x2E80,0x%h_0x%h\n0x2EA0,0x%h_0x%h\n0x2EC0,0x%h_0x%h\n0x2EE0,0x%h_0x%h\n0x2F00,0x%h_0x%h\n0x2F20,0x%h_0x%h\n0x2F40,0x%h_0x%h\n0x2F60,0x%h_0x%h\n0x2F80,0x%h_0x%h\n0x2FA0,0x%h_0x%h\n0x2FC0,0x%h_0x%h\n0x2FE0,0x%h_0x%h\n0x3000,0x%h_0x%h\n0x3020,0x%h_0x%h\n0x3040,0x%h_0x%h\n0x3060,0x%h_0x%h\n0x3080,0x%h_0x%h\n0x30A0,0x%h_0x%h\n0x30C0,0x%h_0x%h\n0x30E0,0x%h_0x%h\n0x3100,0x%h_0x%h\n0x3120,0x%h_0x%h\n0x3140,0x%h_0x%h\n0x3160,0x%h_0x%h\n0x3180,0x%h_0x%h\n0x31A0,0x%h_0x%h\n0x31C0,0x%h_0x%h\n0x31E0,0x%h_0x%h\n0x3200,0x%h_0x%h\n0x3220,0x%h_0x%h\n0x3240,0x%h_0x%h\n0x3260,0x%h_0x%h\n0x3280,0x%h_0x%h\n0x32A0,0x%h_0x%h\n0x32C0,0x%h_0x%h\n0x32E0,0x%h_0x%h\n0x3300,0x%h_0x%h\n0x3320,0x%h_0x%h\n0x3340,0x%h_0x%h\n0x3360,0x%h_0x%h\n0x3380,0x%h_0x%h\n0x33A0,0x%h_0x%h\n0x33C0,0x%h_0x%h\n0x33E0,0x%h_0x%h\n0x3400,0x%h_0x%h\n0x3420,0x%h_0x%h\n0x3440,0x%h_0x%h\n0x3460,0x%h_0x%h\n0x3480,0x%h_0x%h\n0x34A0,0x%h_0x%h\n0x34C0,0x%h_0x%h\n0x34E0,0x%h_0x%h\n0x3500,0x%h_0x%h\n0x3520,0x%h_0x%h\n0x3540,0x%h_0x%h\n0x3560,0x%h_0x%h\n0x3580,0x%h_0x%h\n0x35A0,0x%h_0x%h\n0x35C0,0x%h_0x%h\n0x35E0,0x%h_0x%h\n0x3600,0x%h_0x%h\n0x3620,0x%h_0x%h\n0x3640,0x%h_0x%h\n0x3660,0x%h_0x%h\n0x3680,0x%h_0x%h\n0x36A0,0x%h_0x%h\n0x36C0,0x%h_0x%h\n0x36E0,0x%h_0x%h\n0x3700,0x%h_0x%h\n0x3720,0x%h_0x%h\n0x3740,0x%h_0x%h\n0x3760,0x%h_0x%h\n0x3780,0x%h_0x%h\n0x37A0,0x%h_0x%h\n0x37C0,0x%h_0x%h\n0x37E0,0x%h_0x%h\n0x3800,0x%h_0x%h\n0x3820,0x%h_0x%h\n0x3840,0x%h_0x%h\n0x3860,0x%h_0x%h\n0x3880,0x%h_0x%h\n0x38A0,0x%h_0x%h\n0x38C0,0x%h_0x%h\n0x38E0,0x%h_0x%h\n0x3900,0x%h_0x%h\n0x3920,0x%h_0x%h\n0x3940,0x%h_0x%h\n0x3960,0x%h_0x%h\n0x3980,0x%h_0x%h\n0x39A0,0x%h_0x%h\n0x39C0,0x%h_0x%h\n0x39E0,0x%h_0x%h\n0x3A00,0x%h_0x%h\n0x3A20,0x%h_0x%h\n0x3A40,0x%h_0x%h\n0x3A60,0x%h_0x%h\n0x3A80,0x%h_0x%h\n0x3AA0,0x%h_0x%h\n0x3AC0,0x%h_0x%h\n0x3AE0,0x%h_0x%h\n0x3B00,0x%h_0x%h\n0x3B20,0x%h_0x%h\n0x3B40,0x%h_0x%h\n0x3B60,0x%h_0x%h\n0x3B80,0x%h_0x%h\n0x3BA0,0x%h_0x%h\n0x3BC0,0x%h_0x%h\n0x3BE0,0x%h_0x%h\n0x3C00,0x%h_0x%h\n0x3C20,0x%h_0x%h\n0x3C40,0x%h_0x%h\n0x3C60,0x%h_0x%h\n0x3C80,0x%h_0x%h\n0x3CA0,0x%h_0x%h\n0x3CC0,0x%h_0x%h\n0x3CE0,0x%h_0x%h\n0x3D00,0x%h_0x%h\n0x3D20,0x%h_0x%h\n0x3D40,0x%h_0x%h\n0x3D60,0x%h_0x%h\n0x3D80,0x%h_0x%h\n0x3DA0,0x%h_0x%h\n0x3DC0,0x%h_0x%h\n0x3DE0,0x%h_0x%h\n0x3E00,0x%h_0x%h\n0x3E20,0x%h_0x%h\n0x3E40,0x%h_0x%h\n0x3E60,0x%h_0x%h\n0x3E80,0x%h_0x%h\n0x3EA0,0x%h_0x%h\n0x3EC0,0x%h_0x%h\n0x3EE0,0x%h_0x%h\n0x3F00,0x%h_0x%h\n0x3F20,0x%h_0x%h\n0x3F40,0x%h_0x%h\n0x3F60,0x%h_0x%h\n0x3F80,0x%h_0x%h\n0x3FA0,0x%h_0x%h\n0x3FC0,0x%h_0x%h\n0x3FE0,0x%h_0x%h\n0x4000,0x%h_0x%h\n0x4020,0x%h_0x%h\n0x4040,0x%h_0x%h\n0x4060,0x%h_0x%h\n0x4080,0x%h_0x%h\n0x40A0,0x%h_0x%h\n0x40C0,0x%h_0x%h\n0x40E0,0x%h_0x%h\n0x4100,0x%h_0x%h\n0x4120,0x%h_0x%h\n0x4140,0x%h_0x%h\n0x4160,0x%h_0x%h\n0x4180,0x%h_0x%h\n0x41A0,0x%h_0x%h\n0x41C0,0x%h_0x%h\n0x41E0,0x%h_0x%h\n0x4200,0x%h_0x%h\n0x4220,0x%h_0x%h\n0x4240,0x%h_0x%h\n0x4260,0x%h_0x%h\n0x4280,0x%h_0x%h\n0x42A0,0x%h_0x%h\n0x42C0,0x%h_0x%h\n0x42E0,0x%h_0x%h\n0x4300,0x%h_0x%h\n0x4320,0x%h_0x%h\n0x4340,0x%h_0x%h\n0x4360,0x%h_0x%h\n0x4380,0x%h_0x%h\n0x43A0,0x%h_0x%h\n0x43C0,0x%h_0x%h\n0x43E0,0x%h_0x%h\n0x4400,0x%h_0x%h\n0x4420,0x%h_0x%h\n0x4440,0x%h_0x%h\n0x4460,0x%h_0x%h\n0x4480,0x%h_0x%h\n0x44A0,0x%h_0x%h\n0x44C0,0x%h_0x%h\n0x44E0,0x%h_0x%h\n0x4500,0x%h_0x%h\n0x4520,0x%h_0x%h\n0x4540,0x%h_0x%h\n0x4560,0x%h_0x%h\n0x4580,0x%h_0x%h\n0x45A0,0x%h_0x%h\n0x45C0,0x%h_0x%h\n0x45E0,0x%h_0x%h\n0x4600,0x%h_0x%h\n0x4620,0x%h_0x%h\n0x4640,0x%h_0x%h\n0x4660,0x%h_0x%h\n0x4680,0x%h_0x%h\n0x46A0,0x%h_0x%h\n0x46C0,0x%h_0x%h\n0x46E0,0x%h_0x%h\n0x4700,0x%h_0x%h\n0x4720,0x%h_0x%h\n0x4740,0x%h_0x%h\n0x4760,0x%h_0x%h\n0x4780,0x%h_0x%h\n0x47A0,0x%h_0x%h\n0x47C0,0x%h_0x%h\n0x47E0,0x%h_0x%h\n0x4800,0x%h_0x%h\n0x4820,0x%h_0x%h\n0x4840,0x%h_0x%h\n0x4860,0x%h_0x%h\n0x4880,0x%h_0x%h\n0x48A0,0x%h_0x%h\n0x48C0,0x%h_0x%h\n0x48E0,0x%h_0x%h\n0x4900,0x%h_0x%h\n0x4920,0x%h_0x%h\n0x4940,0x%h_0x%h\n0x4960,0x%h_0x%h\n0x4980,0x%h_0x%h\n0x49A0,0x%h_0x%h\n0x49C0,0x%h_0x%h\n0x49E0,0x%h_0x%h\n0x4A00,0x%h_0x%h\n0x4A20,0x%h_0x%h\n0x4A40,0x%h_0x%h\n0x4A60,0x%h_0x%h\n0x4A80,0x%h_0x%h\n0x4AA0,0x%h_0x%h\n0x4AC0,0x%h_0x%h\n0x4AE0,0x%h_0x%h\n0x4B00,0x%h_0x%h\n0x4B20,0x%h_0x%h\n0x4B40,0x%h_0x%h\n0x4B60,0x%h_0x%h\n0x4B80,0x%h_0x%h\n0x4BA0,0x%h_0x%h\n0x4BC0,0x%h_0x%h\n0x4BE0,0x%h_0x%h\n0x4C00,0x%h_0x%h\n0x4C20,0x%h_0x%h\n0x4C40,0x%h_0x%h\n0x4C60,0x%h_0x%h\n0x4C80,0x%h_0x%h\n0x4CA0,0x%h_0x%h\n0x4CC0,0x%h_0x%h\n0x4CE0,0x%h_0x%h\n0x4D00,0x%h_0x%h\n0x4D20,0x%h_0x%h\n0x4D40,0x%h_0x%h\n0x4D60,0x%h_0x%h\n0x4D80,0x%h_0x%h\n0x4DA0,0x%h_0x%h\n0x4DC0,0x%h_0x%h\n0x4DE0,0x%h_0x%h\n0x4E00,0x%h_0x%h\n0x4E20,0x%h_0x%h\n0x4E40,0x%h_0x%h\n0x4E60,0x%h_0x%h\n0x4E80,0x%h_0x%h\n0x4EA0,0x%h_0x%h\n0x4EC0,0x%h_0x%h\n0x4EE0,0x%h_0x%h\n0x4F00,0x%h_0x%h\n0x4F20,0x%h_0x%h\n0x4F40,0x%h_0x%h\n0x4F60,0x%h_0x%h\n0x4F80,0x%h_0x%h\n0x4FA0,0x%h_0x%h\n0x4FC0,0x%h_0x%h\n0x4FE0,0x%h_0x%h\n0x5000,0x%h_0x%h\n0x5020,0x%h_0x%h\n0x5040,0x%h_0x%h\n0x5060,0x%h_0x%h\n0x5080,0x%h_0x%h\n0x50A0,0x%h_0x%h\n0x50C0,0x%h_0x%h\n0x50E0,0x%h_0x%h\n0x5100,0x%h_0x%h\n0x5120,0x%h_0x%h\n0x5140,0x%h_0x%h\n0x5160,0x%h_0x%h\n0x5180,0x%h_0x%h\n0x51A0,0x%h_0x%h\n0x51C0,0x%h_0x%h\n0x51E0,0x%h_0x%h\n0x5200,0x%h_0x%h\n0x5220,0x%h_0x%h\n0x5240,0x%h_0x%h\n0x5260,0x%h_0x%h\n0x5280,0x%h_0x%h\n0x52A0,0x%h_0x%h\n0x52C0,0x%h_0x%h\n0x52E0,0x%h_0x%h\n0x5300,0x%h_0x%h\n0x5320,0x%h_0x%h\n0x5340,0x%h_0x%h\n0x5360,0x%h_0x%h\n0x5380,0x%h_0x%h\n0x53A0,0x%h_0x%h\n0x53C0,0x%h_0x%h\n0x53E0,0x%h_0x%h\n0x5400,0x%h_0x%h\n0x5420,0x%h_0x%h\n0x5440,0x%h_0x%h\n0x5460,0x%h_0x%h\n0x5480,0x%h_0x%h\n0x54A0,0x%h_0x%h\n0x54C0,0x%h_0x%h\n0x54E0,0x%h_0x%h\n0x5500,0x%h_0x%h\n0x5520,0x%h_0x%h\n0x5540,0x%h_0x%h\n0x5560,0x%h_0x%h\n0x5580,0x%h_0x%h\n0x55A0,0x%h_0x%h\n0x55C0,0x%h_0x%h\n0x55E0,0x%h_0x%h\n0x5600,0x%h_0x%h\n0x5620,0x%h_0x%h\n0x5640,0x%h_0x%h\n0x5660,0x%h_0x%h\n0x5680,0x%h_0x%h\n0x56A0,0x%h_0x%h\n0x56C0,0x%h_0x%h\n0x56E0,0x%h_0x%h\n0x5700,0x%h_0x%h\n0x5720,0x%h_0x%h\n0x5740,0x%h_0x%h\n0x5760,0x%h_0x%h\n0x5780,0x%h_0x%h\n0x57A0,0x%h_0x%h\n0x57C0,0x%h_0x%h\n0x57E0,0x%h_0x%h\n0x5800,0x%h_0x%h\n0x5820,0x%h_0x%h\n0x5840,0x%h_0x%h\n0x5860,0x%h_0x%h\n0x5880,0x%h_0x%h\n0x58A0,0x%h_0x%h\n0x58C0,0x%h_0x%h\n0x58E0,0x%h_0x%h\n0x5900,0x%h_0x%h\n0x5920,0x%h_0x%h\n0x5940,0x%h_0x%h\n0x5960,0x%h_0x%h\n0x5980,0x%h_0x%h\n0x59A0,0x%h_0x%h\n0x59C0,0x%h_0x%h\n0x59E0,0x%h_0x%h\n0x5A00,0x%h_0x%h\n0x5A20,0x%h_0x%h\n0x5A40,0x%h_0x%h\n0x5A60,0x%h_0x%h\n0x5A80,0x%h_0x%h\n0x5AA0,0x%h_0x%h\n0x5AC0,0x%h_0x%h\n0x5AE0,0x%h_0x%h\n0x5B00,0x%h_0x%h\n0x5B20,0x%h_0x%h\n0x5B40,0x%h_0x%h\n0x5B60,0x%h_0x%h\n0x5B80,0x%h_0x%h\n0x5BA0,0x%h_0x%h\n0x5BC0,0x%h_0x%h\n0x5BE0,0x%h_0x%h\n0x5C00,0x%h_0x%h\n0x5C20,0x%h_0x%h\n0x5C40,0x%h_0x%h\n0x5C60,0x%h_0x%h\n0x5C80,0x%h_0x%h\n0x5CA0,0x%h_0x%h\n0x5CC0,0x%h_0x%h\n0x5CE0,0x%h_0x%h\n0x5D00,0x%h_0x%h\n0x5D20,0x%h_0x%h\n0x5D40,0x%h_0x%h\n0x5D60,0x%h_0x%h\n0x5D80,0x%h_0x%h\n0x5DA0,0x%h_0x%h\n0x5DC0,0x%h_0x%h\n0x5DE0,0x%h_0x%h\n0x5E00,0x%h_0x%h\n0x5E20,0x%h_0x%h\n0x5E40,0x%h_0x%h\n0x5E60,0x%h_0x%h\n0x5E80,0x%h_0x%h\n0x5EA0,0x%h_0x%h\n0x5EC0,0x%h_0x%h\n0x5EE0,0x%h_0x%h\n0x5F00,0x%h_0x%h\n0x5F20,0x%h_0x%h\n0x5F40,0x%h_0x%h\n0x5F60,0x%h_0x%h\n0x5F80,0x%h_0x%h\n0x5FA0,0x%h_0x%h\n0x5FC0,0x%h_0x%h\n0x5FE0,0x%h_0x%h\n0x6000,0x%h_0x%h\n0x6020,0x%h_0x%h\n0x6040,0x%h_0x%h\n0x6060,0x%h_0x%h\n0x6080,0x%h_0x%h\n0x60A0,0x%h_0x%h\n0x60C0,0x%h_0x%h\n0x60E0,0x%h_0x%h\n0x6100,0x%h_0x%h\n0x6120,0x%h_0x%h\n0x6140,0x%h_0x%h\n0x6160,0x%h_0x%h\n0x6180,0x%h_0x%h\n0x61A0,0x%h_0x%h\n0x61C0,0x%h_0x%h\n0x61E0,0x%h_0x%h\n0x6200,0x%h_0x%h\n0x6220,0x%h_0x%h\n0x6240,0x%h_0x%h\n0x6260,0x%h_0x%h\n0x6280,0x%h_0x%h\n0x62A0,0x%h_0x%h\n0x62C0,0x%h_0x%h\n0x62E0,0x%h_0x%h\n0x6300,0x%h_0x%h\n0x6320,0x%h_0x%h\n0x6340,0x%h_0x%h\n0x6360,0x%h_0x%h\n0x6380,0x%h_0x%h\n0x63A0,0x%h_0x%h\n0x63C0,0x%h_0x%h\n0x63E0,0x%h_0x%h\n0x6400,0x%h_0x%h\n0x6420,0x%h_0x%h\n0x6440,0x%h_0x%h\n0x6460,0x%h_0x%h\n0x6480,0x%h_0x%h\n0x64A0,0x%h_0x%h\n0x64C0,0x%h_0x%h\n0x64E0,0x%h_0x%h\n0x6500,0x%h_0x%h\n0x6520,0x%h_0x%h\n0x6540,0x%h_0x%h\n0x6560,0x%h_0x%h\n0x6580,0x%h_0x%h\n0x65A0,0x%h_0x%h\n0x65C0,0x%h_0x%h\n0x65E0,0x%h_0x%h\n0x6600,0x%h_0x%h\n0x6620,0x%h_0x%h\n0x6640,0x%h_0x%h\n0x6660,0x%h_0x%h\n0x6680,0x%h_0x%h\n0x66A0,0x%h_0x%h\n0x66C0,0x%h_0x%h\n0x66E0,0x%h_0x%h\n0x6700,0x%h_0x%h\n0x6720,0x%h_0x%h\n0x6740,0x%h_0x%h\n0x6760,0x%h_0x%h\n0x6780,0x%h_0x%h\n0x67A0,0x%h_0x%h\n0x67C0,0x%h_0x%h\n0x67E0,0x%h_0x%h\n0x6800,0x%h_0x%h\n0x6820,0x%h_0x%h\n0x6840,0x%h_0x%h\n0x6860,0x%h_0x%h\n0x6880,0x%h_0x%h\n0x68A0,0x%h_0x%h\n0x68C0,0x%h_0x%h\n0x68E0,0x%h_0x%h\n0x6900,0x%h_0x%h\n0x6920,0x%h_0x%h\n0x6940,0x%h_0x%h\n0x6960,0x%h_0x%h\n0x6980,0x%h_0x%h\n0x69A0,0x%h_0x%h\n0x69C0,0x%h_0x%h\n0x69E0,0x%h_0x%h\n0x6A00,0x%h_0x%h\n0x6A20,0x%h_0x%h\n0x6A40,0x%h_0x%h\n0x6A60,0x%h_0x%h\n0x6A80,0x%h_0x%h\n0x6AA0,0x%h_0x%h\n0x6AC0,0x%h_0x%h\n0x6AE0,0x%h_0x%h\n0x6B00,0x%h_0x%h\n0x6B20,0x%h_0x%h\n0x6B40,0x%h_0x%h\n0x6B60,0x%h_0x%h\n0x6B80,0x%h_0x%h\n0x6BA0,0x%h_0x%h\n0x6BC0,0x%h_0x%h\n0x6BE0,0x%h_0x%h\n0x6C00,0x%h_0x%h\n0x6C20,0x%h_0x%h\n0x6C40,0x%h_0x%h\n0x6C60,0x%h_0x%h\n0x6C80,0x%h_0x%h\n0x6CA0,0x%h_0x%h\n0x6CC0,0x%h_0x%h\n0x6CE0,0x%h_0x%h\n0x6D00,0x%h_0x%h\n0x6D20,0x%h_0x%h\n0x6D40,0x%h_0x%h\n0x6D60,0x%h_0x%h\n0x6D80,0x%h_0x%h\n0x6DA0,0x%h_0x%h\n0x6DC0,0x%h_0x%h\n0x6DE0,0x%h_0x%h\n0x6E00,0x%h_0x%h\n0x6E20,0x%h_0x%h\n0x6E40,0x%h_0x%h\n0x6E60,0x%h_0x%h\n0x6E80,0x%h_0x%h\n0x6EA0,0x%h_0x%h\n0x6EC0,0x%h_0x%h\n0x6EE0,0x%h_0x%h\n0x6F00,0x%h_0x%h\n0x6F20,0x%h_0x%h\n0x6F40,0x%h_0x%h\n0x6F60,0x%h_0x%h\n0x6F80,0x%h_0x%h\n0x6FA0,0x%h_0x%h\n0x6FC0,0x%h_0x%h\n0x6FE0,0x%h_0x%h\n0x7000,0x%h_0x%h\n0x7020,0x%h_0x%h\n0x7040,0x%h_0x%h\n0x7060,0x%h_0x%h\n0x7080,0x%h_0x%h\n0x70A0,0x%h_0x%h\n0x70C0,0x%h_0x%h\n0x70E0,0x%h_0x%h\n0x7100,0x%h_0x%h\n0x7120,0x%h_0x%h\n0x7140,0x%h_0x%h\n0x7160,0x%h_0x%h\n0x7180,0x%h_0x%h\n0x71A0,0x%h_0x%h\n0x71C0,0x%h_0x%h\n0x71E0,0x%h_0x%h\n0x7200,0x%h_0x%h\n0x7220,0x%h_0x%h\n0x7240,0x%h_0x%h\n0x7260,0x%h_0x%h\n0x7280,0x%h_0x%h\n0x72A0,0x%h_0x%h\n0x72C0,0x%h_0x%h\n0x72E0,0x%h_0x%h\n0x7300,0x%h_0x%h\n0x7320,0x%h_0x%h\n0x7340,0x%h_0x%h\n0x7360,0x%h_0x%h\n0x7380,0x%h_0x%h\n0x73A0,0x%h_0x%h\n0x73C0,0x%h_0x%h\n0x73E0,0x%h_0x%h\n0x7400,0x%h_0x%h\n0x7420,0x%h_0x%h\n0x7440,0x%h_0x%h\n0x7460,0x%h_0x%h\n0x7480,0x%h_0x%h\n0x74A0,0x%h_0x%h\n0x74C0,0x%h_0x%h\n0x74E0,0x%h_0x%h\n0x7500,0x%h_0x%h\n0x7520,0x%h_0x%h\n0x7540,0x%h_0x%h\n0x7560,0x%h_0x%h\n0x7580,0x%h_0x%h\n0x75A0,0x%h_0x%h\n0x75C0,0x%h_0x%h\n0x75E0,0x%h_0x%h\n0x7600,0x%h_0x%h\n0x7620,0x%h_0x%h\n0x7640,0x%h_0x%h\n0x7660,0x%h_0x%h\n0x7680,0x%h_0x%h\n0x76A0,0x%h_0x%h\n0x76C0,0x%h_0x%h\n0x76E0,0x%h_0x%h\n0x7700,0x%h_0x%h\n0x7720,0x%h_0x%h\n0x7740,0x%h_0x%h\n0x7760,0x%h_0x%h\n0x7780,0x%h_0x%h\n0x77A0,0x%h_0x%h\n0x77C0,0x%h_0x%h\n0x77E0,0x%h_0x%h\n0x7800,0x%h_0x%h\n0x7820,0x%h_0x%h\n0x7840,0x%h_0x%h\n0x7860,0x%h_0x%h\n0x7880,0x%h_0x%h\n0x78A0,0x%h_0x%h\n0x78C0,0x%h_0x%h\n0x78E0,0x%h_0x%h\n0x7900,0x%h_0x%h\n0x7920,0x%h_0x%h\n0x7940,0x%h_0x%h\n0x7960,0x%h_0x%h\n0x7980,0x%h_0x%h\n0x79A0,0x%h_0x%h\n0x79C0,0x%h_0x%h\n0x79E0,0x%h_0x%h\n0x7A00,0x%h_0x%h\n0x7A20,0x%h_0x%h\n0x7A40,0x%h_0x%h\n0x7A60,0x%h_0x%h\n0x7A80,0x%h_0x%h\n0x7AA0,0x%h_0x%h\n0x7AC0,0x%h_0x%h\n0x7AE0,0x%h_0x%h\n0x7B00,0x%h_0x%h\n0x7B20,0x%h_0x%h\n0x7B40,0x%h_0x%h\n0x7B60,0x%h_0x%h\n0x7B80,0x%h_0x%h\n0x7BA0,0x%h_0x%h\n0x7BC0,0x%h_0x%h\n0x7BE0,0x%h_0x%h\n0x7C00,0x%h_0x%h\n0x7C20,0x%h_0x%h\n0x7C40,0x%h_0x%h\n0x7C60,0x%h_0x%h\n0x7C80,0x%h_0x%h\n0x7CA0,0x%h_0x%h\n0x7CC0,0x%h_0x%h\n0x7CE0,0x%h_0x%h\n0x7D00,0x%h_0x%h\n0x7D20,0x%h_0x%h\n0x7D40,0x%h_0x%h\n0x7D60,0x%h_0x%h\n0x7D80,0x%h_0x%h\n0x7DA0,0x%h_0x%h\n0x7DC0,0x%h_0x%h\n0x7DE0,0x%h_0x%h\n0x7E00,0x%h_0x%h\n0x7E20,0x%h_0x%h\n0x7E40,0x%h_0x%h\n0x7E60,0x%h_0x%h\n0x7E80,0x%h_0x%h\n0x7EA0,0x%h_0x%h\n0x7EC0,0x%h_0x%h\n0x7EE0,0x%h_0x%h\n0x7F00,0x%h_0x%h\n0x7F20,0x%h_0x%h\n0x7F40,0x%h_0x%h\n0x7F60,0x%h_0x%h\n0x7F80,0x%h_0x%h\n0x7FA0,0x%h_0x%h\n0x7FC0,0x%h_0x%h\n0x7FE0,0x%h_0x%h\n0x8000,0x%h_0x%h\n0x8020,0x%h_0x%h\n0x8040,0x%h_0x%h\n0x8060,0x%h_0x%h\n0x8080,0x%h_0x%h\n0x80A0,0x%h_0x%h\n0x80C0,0x%h_0x%h\n0x80E0,0x%h_0x%h\n0x8100,0x%h_0x%h\n0x8120,0x%h_0x%h\n0x8140,0x%h_0x%h\n0x8160,0x%h_0x%h\n0x8180,0x%h_0x%h\n0x81A0,0x%h_0x%h\n0x81C0,0x%h_0x%h\n0x81E0,0x%h_0x%h\n0x8200,0x%h_0x%h\n0x8220,0x%h_0x%h\n0x8240,0x%h_0x%h\n0x8260,0x%h_0x%h\n0x8280,0x%h_0x%h\n0x82A0,0x%h_0x%h\n0x82C0,0x%h_0x%h\n0x82E0,0x%h_0x%h\n0x8300,0x%h_0x%h\n0x8320,0x%h_0x%h\n0x8340,0x%h_0x%h\n0x8360,0x%h_0x%h\n0x8380,0x%h_0x%h\n0x83A0,0x%h_0x%h\n0x83C0,0x%h_0x%h\n0x83E0,0x%h_0x%h\n0x8400,0x%h_0x%h\n0x8420,0x%h_0x%h\n0x8440,0x%h_0x%h\n0x8460,0x%h_0x%h\n0x8480,0x%h_0x%h\n0x84A0,0x%h_0x%h\n0x84C0,0x%h_0x%h\n0x84E0,0x%h_0x%h\n0x8500,0x%h_0x%h\n0x8520,0x%h_0x%h\n0x8540,0x%h_0x%h\n0x8560,0x%h_0x%h\n0x8580,0x%h_0x%h\n0x85A0,0x%h_0x%h\n0x85C0,0x%h_0x%h\n0x85E0,0x%h_0x%h\n0x8600,0x%h_0x%h\n0x8620,0x%h_0x%h\n0x8640,0x%h_0x%h\n0x8660,0x%h_0x%h\n0x8680,0x%h_0x%h\n0x86A0,0x%h_0x%h\n0x86C0,0x%h_0x%h\n0x86E0,0x%h_0x%h\n0x8700,0x%h_0x%h\n0x8720,0x%h_0x%h\n0x8740,0x%h_0x%h\n0x8760,0x%h_0x%h\n0x8780,0x%h_0x%h\n0x87A0,0x%h_0x%h\n0x87C0,0x%h_0x%h\n0x87E0,0x%h_0x%h\n0x8800,0x%h_0x%h\n0x8820,0x%h_0x%h\n0x8840,0x%h_0x%h\n0x8860,0x%h_0x%h\n0x8880,0x%h_0x%h\n0x88A0,0x%h_0x%h\n0x88C0,0x%h_0x%h\n0x88E0,0x%h_0x%h\n0x8900,0x%h_0x%h\n0x8920,0x%h_0x%h\n0x8940,0x%h_0x%h\n0x8960,0x%h_0x%h\n0x8980,0x%h_0x%h\n0x89A0,0x%h_0x%h\n0x89C0,0x%h_0x%h\n0x89E0,0x%h_0x%h\n0x8A00,0x%h_0x%h\n0x8A20,0x%h_0x%h\n0x8A40,0x%h_0x%h\n0x8A60,0x%h_0x%h\n0x8A80,0x%h_0x%h\n0x8AA0,0x%h_0x%h\n0x8AC0,0x%h_0x%h\n0x8AE0,0x%h_0x%h\n0x8B00,0x%h_0x%h\n0x8B20,0x%h_0x%h\n0x8B40,0x%h_0x%h\n0x8B60,0x%h_0x%h\n0x8B80,0x%h_0x%h\n0x8BA0,0x%h_0x%h\n0x8BC0,0x%h_0x%h\n0x8BE0,0x%h_0x%h\n0x8C00,0x%h_0x%h\n0x8C20,0x%h_0x%h\n0x8C40,0x%h_0x%h\n0x8C60,0x%h_0x%h\n0x8C80,0x%h_0x%h\n0x8CA0,0x%h_0x%h\n0x8CC0,0x%h_0x%h\n0x8CE0,0x%h_0x%h\n0x8D00,0x%h_0x%h\n0x8D20,0x%h_0x%h\n0x8D40,0x%h_0x%h\n0x8D60,0x%h_0x%h\n0x8D80,0x%h_0x%h\n0x8DA0,0x%h_0x%h\n0x8DC0,0x%h_0x%h\n0x8DE0,0x%h_0x%h\n0x8E00,0x%h_0x%h\n0x8E20,0x%h_0x%h\n0x8E40,0x%h_0x%h\n0x8E60,0x%h_0x%h\n0x8E80,0x%h_0x%h\n0x8EA0,0x%h_0x%h\n0x8EC0,0x%h_0x%h\n0x8EE0,0x%h_0x%h\n0x8F00,0x%h_0x%h\n0x8F20,0x%h_0x%h\n0x8F40,0x%h_0x%h\n0x8F60,0x%h_0x%h\n0x8F80,0x%h_0x%h\n0x8FA0,0x%h_0x%h\n0x8FC0,0x%h_0x%h\n0x8FE0,0x%h_0x%h\n0x9000,0x%h_0x%h\n0x9020,0x%h_0x%h\n0x9040,0x%h_0x%h\n0x9060,0x%h_0x%h\n0x9080,0x%h_0x%h\n0x90A0,0x%h_0x%h\n0x90C0,0x%h_0x%h\n0x90E0,0x%h_0x%h\n0x9100,0x%h_0x%h\n0x9120,0x%h_0x%h\n0x9140,0x%h_0x%h\n0x9160,0x%h_0x%h\n0x9180,0x%h_0x%h\n0x91A0,0x%h_0x%h\n0x91C0,0x%h_0x%h\n0x91E0,0x%h_0x%h\n0x9200,0x%h_0x%h\n0x9220,0x%h_0x%h\n0x9240,0x%h_0x%h\n0x9260,0x%h_0x%h\n0x9280,0x%h_0x%h\n0x92A0,0x%h_0x%h\n0x92C0,0x%h_0x%h\n0x92E0,0x%h_0x%h\n0x9300,0x%h_0x%h\n0x9320,0x%h_0x%h\n0x9340,0x%h_0x%h\n0x9360,0x%h_0x%h\n0x9380,0x%h_0x%h\n0x93A0,0x%h_0x%h\n0x93C0,0x%h_0x%h\n0x93E0,0x%h_0x%h\n0x9400,0x%h_0x%h\n0x9420,0x%h_0x%h\n0x9440,0x%h_0x%h\n0x9460,0x%h_0x%h\n0x9480,0x%h_0x%h\n0x94A0,0x%h_0x%h\n0x94C0,0x%h_0x%h\n0x94E0,0x%h_0x%h\n0x9500,0x%h_0x%h\n0x9520,0x%h_0x%h\n0x9540,0x%h_0x%h\n0x9560,0x%h_0x%h\n0x9580,0x%h_0x%h\n0x95A0,0x%h_0x%h\n0x95C0,0x%h_0x%h\n0x95E0,0x%h_0x%h\n0x9600,0x%h_0x%h\n0x9620,0x%h_0x%h\n0x9640,0x%h_0x%h\n0x9660,0x%h_0x%h\n0x9680,0x%h_0x%h\n0x96A0,0x%h_0x%h\n0x96C0,0x%h_0x%h\n0x96E0,0x%h_0x%h\n0x9700,0x%h_0x%h\n0x9720,0x%h_0x%h\n0x9740,0x%h_0x%h\n0x9760,0x%h_0x%h\n0x9780,0x%h_0x%h\n0x97A0,0x%h_0x%h\n0x97C0,0x%h_0x%h\n0x97E0,0x%h_0x%h\n0x9800,0x%h_0x%h\n0x9820,0x%h_0x%h\n0x9840,0x%h_0x%h\n0x9860,0x%h_0x%h\n0x9880,0x%h_0x%h\n0x98A0,0x%h_0x%h\n0x98C0,0x%h_0x%h\n0x98E0,0x%h_0x%h\n0x9900,0x%h_0x%h\n0x9920,0x%h_0x%h\n0x9940,0x%h_0x%h\n0x9960,0x%h_0x%h\n0x9980,0x%h_0x%h\n0x99A0,0x%h_0x%h\n0x99C0,0x%h_0x%h\n0x99E0,0x%h_0x%h\n0x9A00,0x%h_0x%h\n0x9A20,0x%h_0x%h\n0x9A40,0x%h_0x%h\n0x9A60,0x%h_0x%h\n0x9A80,0x%h_0x%h\n0x9AA0,0x%h_0x%h\n0x9AC0,0x%h_0x%h\n0x9AE0,0x%h_0x%h\n0x9B00,0x%h_0x%h\n0x9B20,0x%h_0x%h\n0x9B40,0x%h_0x%h\n0x9B60,0x%h_0x%h\n0x9B80,0x%h_0x%h\n0x9BA0,0x%h_0x%h\n0x9BC0,0x%h_0x%h\n0x9BE0,0x%h_0x%h\n0x9C00,0x%h_0x%h\n0x9C20,0x%h_0x%h\n0x9C40,0x%h_0x%h\n0x9C60,0x%h_0x%h\n0x9C80,0x%h_0x%h\n0x9CA0,0x%h_0x%h\n0x9CC0,0x%h_0x%h\n0x9CE0,0x%h_0x%h\n0x9D00,0x%h_0x%h\n0x9D20,0x%h_0x%h\n0x9D40,0x%h_0x%h\n0x9D60,0x%h_0x%h\n0x9D80,0x%h_0x%h\n0x9DA0,0x%h_0x%h\n0x9DC0,0x%h_0x%h\n0x9DE0,0x%h_0x%h\n0x9E00,0x%h_0x%h\n0x9E20,0x%h_0x%h\n0x9E40,0x%h_0x%h\n0x9E60,0x%h_0x%h\n0x9E80,0x%h_0x%h\n0x9EA0,0x%h_0x%h\n0x9EC0,0x%h_0x%h\n0x9EE0,0x%h_0x%h\n0x9F00,0x%h_0x%h\n0x9F20,0x%h_0x%h\n0x9F40,0x%h_0x%h\n0x9F60,0x%h_0x%h\n0x9F80,0x%h_0x%h\n0x9FA0,0x%h_0x%h\n0x9FC0,0x%h_0x%h\n0x9FE0,0x%h_0x%h\n0xA000,0x%h_0x%h\n0xA020,0x%h_0x%h\n0xA040,0x%h_0x%h\n0xA060,0x%h_0x%h\n0xA080,0x%h_0x%h\n0xA0A0,0x%h_0x%h\n0xA0C0,0x%h_0x%h\n0xA0E0,0x%h_0x%h\n0xA100,0x%h_0x%h\n0xA120,0x%h_0x%h\n0xA140,0x%h_0x%h\n0xA160,0x%h_0x%h\n0xA180,0x%h_0x%h\n0xA1A0,0x%h_0x%h\n0xA1C0,0x%h_0x%h\n0xA1E0,0x%h_0x%h\n0xA200,0x%h_0x%h\n0xA220,0x%h_0x%h\n0xA240,0x%h_0x%h\n0xA260,0x%h_0x%h\n0xA280,0x%h_0x%h\n0xA2A0,0x%h_0x%h\n0xA2C0,0x%h_0x%h\n0xA2E0,0x%h_0x%h\n0xA300,0x%h_0x%h\n0xA320,0x%h_0x%h\n0xA340,0x%h_0x%h\n0xA360,0x%h_0x%h\n0xA380,0x%h_0x%h\n0xA3A0,0x%h_0x%h\n0xA3C0,0x%h_0x%h\n0xA3E0,0x%h_0x%h\n0xA400,0x%h_0x%h\n0xA420,0x%h_0x%h\n0xA440,0x%h_0x%h\n0xA460,0x%h_0x%h\n0xA480,0x%h_0x%h\n0xA4A0,0x%h_0x%h\n0xA4C0,0x%h_0x%h\n0xA4E0,0x%h_0x%h\n0xA500,0x%h_0x%h\n0xA520,0x%h_0x%h\n0xA540,0x%h_0x%h\n0xA560,0x%h_0x%h\n0xA580,0x%h_0x%h\n0xA5A0,0x%h_0x%h\n0xA5C0,0x%h_0x%h\n0xA5E0,0x%h_0x%h\n0xA600,0x%h_0x%h\n0xA620,0x%h_0x%h\n0xA640,0x%h_0x%h\n0xA660,0x%h_0x%h\n0xA680,0x%h_0x%h\n0xA6A0,0x%h_0x%h\n0xA6C0,0x%h_0x%h\n0xA6E0,0x%h_0x%h\n0xA700,0x%h_0x%h\n0xA720,0x%h_0x%h\n0xA740,0x%h_0x%h\n0xA760,0x%h_0x%h\n0xA780,0x%h_0x%h\n0xA7A0,0x%h_0x%h\n0xA7C0,0x%h_0x%h\n0xA7E0,0x%h_0x%h\n0xA800,0x%h_0x%h\n0xA820,0x%h_0x%h\n0xA840,0x%h_0x%h\n0xA860,0x%h_0x%h\n0xA880,0x%h_0x%h\n0xA8A0,0x%h_0x%h\n0xA8C0,0x%h_0x%h\n0xA8E0,0x%h_0x%h\n0xA900,0x%h_0x%h\n0xA920,0x%h_0x%h\n0xA940,0x%h_0x%h\n0xA960,0x%h_0x%h\n0xA980,0x%h_0x%h\n0xA9A0,0x%h_0x%h\n0xA9C0,0x%h_0x%h\n0xA9E0,0x%h_0x%h\n0xAA00,0x%h_0x%h\n0xAA20,0x%h_0x%h\n0xAA40,0x%h_0x%h\n0xAA60,0x%h_0x%h\n0xAA80,0x%h_0x%h\n0xAAA0,0x%h_0x%h\n0xAAC0,0x%h_0x%h\n0xAAE0,0x%h_0x%h\n0xAB00,0x%h_0x%h\n0xAB20,0x%h_0x%h\n0xAB40,0x%h_0x%h\n0xAB60,0x%h_0x%h\n0xAB80,0x%h_0x%h\n0xABA0,0x%h_0x%h\n0xABC0,0x%h_0x%h\n0xABE0,0x%h_0x%h\n0xAC00,0x%h_0x%h\n0xAC20,0x%h_0x%h\n0xAC40,0x%h_0x%h\n0xAC60,0x%h_0x%h\n0xAC80,0x%h_0x%h\n0xACA0,0x%h_0x%h\n0xACC0,0x%h_0x%h\n0xACE0,0x%h_0x%h\n0xAD00,0x%h_0x%h\n0xAD20,0x%h_0x%h\n0xAD40,0x%h_0x%h\n0xAD60,0x%h_0x%h\n0xAD80,0x%h_0x%h\n0xADA0,0x%h_0x%h\n0xADC0,0x%h_0x%h\n0xADE0,0x%h_0x%h\n0xAE00,0x%h_0x%h\n0xAE20,0x%h_0x%h\n0xAE40,0x%h_0x%h\n0xAE60,0x%h_0x%h\n0xAE80,0x%h_0x%h\n0xAEA0,0x%h_0x%h\n0xAEC0,0x%h_0x%h\n0xAEE0,0x%h_0x%h\n0xAF00,0x%h_0x%h\n0xAF20,0x%h_0x%h\n0xAF40,0x%h_0x%h\n0xAF60,0x%h_0x%h\n0xAF80,0x%h_0x%h\n0xAFA0,0x%h_0x%h\n0xAFC0,0x%h_0x%h\n0xAFE0,0x%h_0x%h\n0xB000,0x%h_0x%h\n0xB020,0x%h_0x%h\n0xB040,0x%h_0x%h\n0xB060,0x%h_0x%h\n0xB080,0x%h_0x%h\n0xB0A0,0x%h_0x%h\n0xB0C0,0x%h_0x%h\n0xB0E0,0x%h_0x%h\n0xB100,0x%h_0x%h\n0xB120,0x%h_0x%h\n0xB140,0x%h_0x%h\n0xB160,0x%h_0x%h\n0xB180,0x%h_0x%h\n0xB1A0,0x%h_0x%h\n0xB1C0,0x%h_0x%h\n0xB1E0,0x%h_0x%h\n0xB200,0x%h_0x%h\n0xB220,0x%h_0x%h\n0xB240,0x%h_0x%h\n0xB260,0x%h_0x%h\n0xB280,0x%h_0x%h\n0xB2A0,0x%h_0x%h\n0xB2C0,0x%h_0x%h\n0xB2E0,0x%h_0x%h\n0xB300,0x%h_0x%h\n0xB320,0x%h_0x%h\n0xB340,0x%h_0x%h\n0xB360,0x%h_0x%h\n0xB380,0x%h_0x%h\n0xB3A0,0x%h_0x%h\n0xB3C0,0x%h_0x%h\n0xB3E0,0x%h_0x%h\n0xB400,0x%h_0x%h\n0xB420,0x%h_0x%h\n0xB440,0x%h_0x%h\n0xB460,0x%h_0x%h\n0xB480,0x%h_0x%h\n0xB4A0,0x%h_0x%h\n0xB4C0,0x%h_0x%h\n0xB4E0,0x%h_0x%h\n0xB500,0x%h_0x%h\n0xB520,0x%h_0x%h\n0xB540,0x%h_0x%h\n0xB560,0x%h_0x%h\n0xB580,0x%h_0x%h\n0xB5A0,0x%h_0x%h\n0xB5C0,0x%h_0x%h\n0xB5E0,0x%h_0x%h\n0xB600,0x%h_0x%h\n0xB620,0x%h_0x%h\n0xB640,0x%h_0x%h\n0xB660,0x%h_0x%h\n0xB680,0x%h_0x%h\n0xB6A0,0x%h_0x%h\n0xB6C0,0x%h_0x%h\n0xB6E0,0x%h_0x%h\n0xB700,0x%h_0x%h\n0xB720,0x%h_0x%h\n0xB740,0x%h_0x%h\n0xB760,0x%h_0x%h\n0xB780,0x%h_0x%h\n0xB7A0,0x%h_0x%h\n0xB7C0,0x%h_0x%h\n0xB7E0,0x%h_0x%h\n0xB800,0x%h_0x%h\n0xB820,0x%h_0x%h\n0xB840,0x%h_0x%h\n0xB860,0x%h_0x%h\n0xB880,0x%h_0x%h\n0xB8A0,0x%h_0x%h\n0xB8C0,0x%h_0x%h\n0xB8E0,0x%h_0x%h\n0xB900,0x%h_0x%h\n0xB920,0x%h_0x%h\n0xB940,0x%h_0x%h\n0xB960,0x%h_0x%h\n0xB980,0x%h_0x%h\n0xB9A0,0x%h_0x%h\n0xB9C0,0x%h_0x%h\n0xB9E0,0x%h_0x%h\n0xBA00,0x%h_0x%h\n0xBA20,0x%h_0x%h\n0xBA40,0x%h_0x%h\n0xBA60,0x%h_0x%h\n0xBA80,0x%h_0x%h\n0xBAA0,0x%h_0x%h\n0xBAC0,0x%h_0x%h\n0xBAE0,0x%h_0x%h\n0xBB00,0x%h_0x%h\n0xBB20,0x%h_0x%h\n0xBB40,0x%h_0x%h\n0xBB60,0x%h_0x%h\n0xBB80,0x%h_0x%h\n0xBBA0,0x%h_0x%h\n0xBBC0,0x%h_0x%h\n0xBBE0,0x%h_0x%h\n0xBC00,0x%h_0x%h\n0xBC20,0x%h_0x%h\n0xBC40,0x%h_0x%h\n0xBC60,0x%h_0x%h\n0xBC80,0x%h_0x%h\n0xBCA0,0x%h_0x%h\n0xBCC0,0x%h_0x%h\n0xBCE0,0x%h_0x%h\n0xBD00,0x%h_0x%h\n0xBD20,0x%h_0x%h\n0xBD40,0x%h_0x%h\n0xBD60,0x%h_0x%h\n0xBD80,0x%h_0x%h\n0xBDA0,0x%h_0x%h\n0xBDC0,0x%h_0x%h\n0xBDE0,0x%h_0x%h\n0xBE00,0x%h_0x%h\n0xBE20,0x%h_0x%h\n0xBE40,0x%h_0x%h\n0xBE60,0x%h_0x%h\n0xBE80,0x%h_0x%h\n0xBEA0,0x%h_0x%h\n0xBEC0,0x%h_0x%h\n0xBEE0,0x%h_0x%h\n0xBF00,0x%h_0x%h\n0xBF20,0x%h_0x%h\n0xBF40,0x%h_0x%h\n0xBF60,0x%h_0x%h\n0xBF80,0x%h_0x%h\n0xBFA0,0x%h_0x%h\n0xBFC0,0x%h_0x%h\n0xBFE0,0x%h_0x%h\n0xC000,0x%h_0x%h\n0xC020,0x%h_0x%h\n0xC040,0x%h_0x%h\n0xC060,0x%h_0x%h\n0xC080,0x%h_0x%h\n0xC0A0,0x%h_0x%h\n0xC0C0,0x%h_0x%h\n0xC0E0,0x%h_0x%h\n0xC100,0x%h_0x%h\n0xC120,0x%h_0x%h\n0xC140,0x%h_0x%h\n0xC160,0x%h_0x%h\n0xC180,0x%h_0x%h\n0xC1A0,0x%h_0x%h\n0xC1C0,0x%h_0x%h\n0xC1E0,0x%h_0x%h\n0xC200,0x%h_0x%h\n0xC220,0x%h_0x%h\n0xC240,0x%h_0x%h\n0xC260,0x%h_0x%h\n0xC280,0x%h_0x%h\n0xC2A0,0x%h_0x%h\n0xC2C0,0x%h_0x%h\n0xC2E0,0x%h_0x%h\n0xC300,0x%h_0x%h\n0xC320,0x%h_0x%h\n0xC340,0x%h_0x%h\n0xC360,0x%h_0x%h\n0xC380,0x%h_0x%h\n0xC3A0,0x%h_0x%h\n0xC3C0,0x%h_0x%h\n0xC3E0,0x%h_0x%h\n0xC400,0x%h_0x%h\n0xC420,0x%h_0x%h\n0xC440,0x%h_0x%h\n0xC460,0x%h_0x%h\n0xC480,0x%h_0x%h\n0xC4A0,0x%h_0x%h\n0xC4C0,0x%h_0x%h\n0xC4E0,0x%h_0x%h\n0xC500,0x%h_0x%h\n0xC520,0x%h_0x%h\n0xC540,0x%h_0x%h\n0xC560,0x%h_0x%h\n0xC580,0x%h_0x%h\n0xC5A0,0x%h_0x%h\n0xC5C0,0x%h_0x%h\n0xC5E0,0x%h_0x%h\n0xC600,0x%h_0x%h\n0xC620,0x%h_0x%h\n0xC640,0x%h_0x%h\n0xC660,0x%h_0x%h\n0xC680,0x%h_0x%h\n0xC6A0,0x%h_0x%h\n0xC6C0,0x%h_0x%h\n0xC6E0,0x%h_0x%h\n0xC700,0x%h_0x%h\n0xC720,0x%h_0x%h\n0xC740,0x%h_0x%h\n0xC760,0x%h_0x%h\n0xC780,0x%h_0x%h\n0xC7A0,0x%h_0x%h\n0xC7C0,0x%h_0x%h\n0xC7E0,0x%h_0x%h\n0xC800,0x%h_0x%h\n0xC820,0x%h_0x%h\n0xC840,0x%h_0x%h\n0xC860,0x%h_0x%h\n0xC880,0x%h_0x%h\n0xC8A0,0x%h_0x%h\n0xC8C0,0x%h_0x%h\n0xC8E0,0x%h_0x%h\n0xC900,0x%h_0x%h\n0xC920,0x%h_0x%h\n0xC940,0x%h_0x%h\n0xC960,0x%h_0x%h\n0xC980,0x%h_0x%h\n0xC9A0,0x%h_0x%h\n0xC9C0,0x%h_0x%h\n0xC9E0,0x%h_0x%h\n0xCA00,0x%h_0x%h\n0xCA20,0x%h_0x%h\n0xCA40,0x%h_0x%h\n0xCA60,0x%h_0x%h\n0xCA80,0x%h_0x%h\n0xCAA0,0x%h_0x%h\n0xCAC0,0x%h_0x%h\n0xCAE0,0x%h_0x%h\n0xCB00,0x%h_0x%h\n0xCB20,0x%h_0x%h\n0xCB40,0x%h_0x%h\n0xCB60,0x%h_0x%h\n0xCB80,0x%h_0x%h\n0xCBA0,0x%h_0x%h\n0xCBC0,0x%h_0x%h\n0xCBE0,0x%h_0x%h\n0xCC00,0x%h_0x%h\n0xCC20,0x%h_0x%h\n0xCC40,0x%h_0x%h\n0xCC60,0x%h_0x%h\n0xCC80,0x%h_0x%h\n0xCCA0,0x%h_0x%h\n0xCCC0,0x%h_0x%h\n0xCCE0,0x%h_0x%h\n0xCD00,0x%h_0x%h\n0xCD20,0x%h_0x%h\n0xCD40,0x%h_0x%h\n0xCD60,0x%h_0x%h\n0xCD80,0x%h_0x%h\n0xCDA0,0x%h_0x%h\n0xCDC0,0x%h_0x%h\n0xCDE0,0x%h_0x%h\n0xCE00,0x%h_0x%h\n0xCE20,0x%h_0x%h\n0xCE40,0x%h_0x%h\n0xCE60,0x%h_0x%h\n0xCE80,0x%h_0x%h\n0xCEA0,0x%h_0x%h\n0xCEC0,0x%h_0x%h\n0xCEE0,0x%h_0x%h\n0xCF00,0x%h_0x%h\n0xCF20,0x%h_0x%h\n0xCF40,0x%h_0x%h\n0xCF60,0x%h_0x%h\n0xCF80,0x%h_0x%h\n0xCFA0,0x%h_0x%h\n0xCFC0,0x%h_0x%h\n0xCFE0,0x%h_0x%h\n0xD000,0x%h_0x%h\n0xD020,0x%h_0x%h\n0xD040,0x%h_0x%h\n0xD060,0x%h_0x%h\n0xD080,0x%h_0x%h\n0xD0A0,0x%h_0x%h\n0xD0C0,0x%h_0x%h\n0xD0E0,0x%h_0x%h\n0xD100,0x%h_0x%h\n0xD120,0x%h_0x%h\n0xD140,0x%h_0x%h\n0xD160,0x%h_0x%h\n0xD180,0x%h_0x%h\n0xD1A0,0x%h_0x%h\n0xD1C0,0x%h_0x%h\n0xD1E0,0x%h_0x%h\n0xD200,0x%h_0x%h\n0xD220,0x%h_0x%h\n0xD240,0x%h_0x%h\n0xD260,0x%h_0x%h\n0xD280,0x%h_0x%h\n0xD2A0,0x%h_0x%h\n0xD2C0,0x%h_0x%h\n0xD2E0,0x%h_0x%h\n0xD300,0x%h_0x%h\n0xD320,0x%h_0x%h\n0xD340,0x%h_0x%h\n0xD360,0x%h_0x%h\n0xD380,0x%h_0x%h\n0xD3A0,0x%h_0x%h\n0xD3C0,0x%h_0x%h\n0xD3E0,0x%h_0x%h\n0xD400,0x%h_0x%h\n0xD420,0x%h_0x%h\n0xD440,0x%h_0x%h\n0xD460,0x%h_0x%h\n0xD480,0x%h_0x%h\n0xD4A0,0x%h_0x%h\n0xD4C0,0x%h_0x%h\n0xD4E0,0x%h_0x%h\n0xD500,0x%h_0x%h\n0xD520,0x%h_0x%h\n0xD540,0x%h_0x%h\n0xD560,0x%h_0x%h\n0xD580,0x%h_0x%h\n0xD5A0,0x%h_0x%h\n0xD5C0,0x%h_0x%h\n0xD5E0,0x%h_0x%h\n0xD600,0x%h_0x%h\n0xD620,0x%h_0x%h\n0xD640,0x%h_0x%h\n0xD660,0x%h_0x%h\n0xD680,0x%h_0x%h\n0xD6A0,0x%h_0x%h\n0xD6C0,0x%h_0x%h\n0xD6E0,0x%h_0x%h\n0xD700,0x%h_0x%h\n0xD720,0x%h_0x%h\n0xD740,0x%h_0x%h\n0xD760,0x%h_0x%h\n0xD780,0x%h_0x%h\n0xD7A0,0x%h_0x%h\n0xD7C0,0x%h_0x%h\n0xD7E0,0x%h_0x%h\n0xD800,0x%h_0x%h\n0xD820,0x%h_0x%h\n0xD840,0x%h_0x%h\n0xD860,0x%h_0x%h\n0xD880,0x%h_0x%h\n0xD8A0,0x%h_0x%h\n0xD8C0,0x%h_0x%h\n0xD8E0,0x%h_0x%h\n0xD900,0x%h_0x%h\n0xD920,0x%h_0x%h\n0xD940,0x%h_0x%h\n0xD960,0x%h_0x%h\n0xD980,0x%h_0x%h\n0xD9A0,0x%h_0x%h\n0xD9C0,0x%h_0x%h\n0xD9E0,0x%h_0x%h\n0xDA00,0x%h_0x%h\n0xDA20,0x%h_0x%h\n0xDA40,0x%h_0x%h\n0xDA60,0x%h_0x%h\n0xDA80,0x%h_0x%h\n0xDAA0,0x%h_0x%h\n0xDAC0,0x%h_0x%h\n0xDAE0,0x%h_0x%h\n0xDB00,0x%h_0x%h\n0xDB20,0x%h_0x%h\n0xDB40,0x%h_0x%h\n0xDB60,0x%h_0x%h\n0xDB80,0x%h_0x%h\n0xDBA0,0x%h_0x%h\n0xDBC0,0x%h_0x%h\n0xDBE0,0x%h_0x%h\n0xDC00,0x%h_0x%h\n0xDC20,0x%h_0x%h\n0xDC40,0x%h_0x%h\n0xDC60,0x%h_0x%h\n0xDC80,0x%h_0x%h\n0xDCA0,0x%h_0x%h\n0xDCC0,0x%h_0x%h\n0xDCE0,0x%h_0x%h\n0xDD00,0x%h_0x%h\n0xDD20,0x%h_0x%h\n0xDD40,0x%h_0x%h\n0xDD60,0x%h_0x%h\n0xDD80,0x%h_0x%h\n0xDDA0,0x%h_0x%h\n0xDDC0,0x%h_0x%h\n0xDDE0,0x%h_0x%h\n0xDE00,0x%h_0x%h\n0xDE20,0x%h_0x%h\n0xDE40,0x%h_0x%h\n0xDE60,0x%h_0x%h\n0xDE80,0x%h_0x%h\n0xDEA0,0x%h_0x%h\n0xDEC0,0x%h_0x%h\n0xDEE0,0x%h_0x%h\n0xDF00,0x%h_0x%h\n0xDF20,0x%h_0x%h\n0xDF40,0x%h_0x%h\n0xDF60,0x%h_0x%h\n0xDF80,0x%h_0x%h\n0xDFA0,0x%h_0x%h\n0xDFC0,0x%h_0x%h\n0xDFE0,0x%h_0x%h\n0xE000,0x%h_0x%h\n0xE020,0x%h_0x%h\n0xE040,0x%h_0x%h\n0xE060,0x%h_0x%h\n0xE080,0x%h_0x%h\n0xE0A0,0x%h_0x%h\n0xE0C0,0x%h_0x%h\n0xE0E0,0x%h_0x%h\n0xE100,0x%h_0x%h\n0xE120,0x%h_0x%h\n0xE140,0x%h_0x%h\n0xE160,0x%h_0x%h\n0xE180,0x%h_0x%h\n0xE1A0,0x%h_0x%h\n0xE1C0,0x%h_0x%h\n0xE1E0,0x%h_0x%h\n0xE200,0x%h_0x%h\n0xE220,0x%h_0x%h\n0xE240,0x%h_0x%h\n0xE260,0x%h_0x%h\n0xE280,0x%h_0x%h\n0xE2A0,0x%h_0x%h\n0xE2C0,0x%h_0x%h\n0xE2E0,0x%h_0x%h\n0xE300,0x%h_0x%h\n0xE320,0x%h_0x%h\n0xE340,0x%h_0x%h\n0xE360,0x%h_0x%h\n0xE380,0x%h_0x%h\n0xE3A0,0x%h_0x%h\n0xE3C0,0x%h_0x%h\n0xE3E0,0x%h_0x%h\n0xE400,0x%h_0x%h\n0xE420,0x%h_0x%h\n0xE440,0x%h_0x%h\n0xE460,0x%h_0x%h\n0xE480,0x%h_0x%h\n0xE4A0,0x%h_0x%h\n0xE4C0,0x%h_0x%h\n0xE4E0,0x%h_0x%h\n0xE500,0x%h_0x%h\n0xE520,0x%h_0x%h\n0xE540,0x%h_0x%h\n0xE560,0x%h_0x%h\n0xE580,0x%h_0x%h\n0xE5A0,0x%h_0x%h\n0xE5C0,0x%h_0x%h\n0xE5E0,0x%h_0x%h\n0xE600,0x%h_0x%h\n0xE620,0x%h_0x%h\n0xE640,0x%h_0x%h\n0xE660,0x%h_0x%h\n0xE680,0x%h_0x%h\n0xE6A0,0x%h_0x%h\n0xE6C0,0x%h_0x%h\n0xE6E0,0x%h_0x%h\n0xE700,0x%h_0x%h\n0xE720,0x%h_0x%h\n0xE740,0x%h_0x%h\n0xE760,0x%h_0x%h\n0xE780,0x%h_0x%h\n0xE7A0,0x%h_0x%h\n0xE7C0,0x%h_0x%h\n0xE7E0,0x%h_0x%h\n0xE800,0x%h_0x%h\n0xE820,0x%h_0x%h\n0xE840,0x%h_0x%h\n0xE860,0x%h_0x%h\n0xE880,0x%h_0x%h\n0xE8A0,0x%h_0x%h\n0xE8C0,0x%h_0x%h\n0xE8E0,0x%h_0x%h\n0xE900,0x%h_0x%h\n0xE920,0x%h_0x%h\n0xE940,0x%h_0x%h\n0xE960,0x%h_0x%h\n0xE980,0x%h_0x%h\n0xE9A0,0x%h_0x%h\n0xE9C0,0x%h_0x%h\n0xE9E0,0x%h_0x%h\n0xEA00,0x%h_0x%h\n0xEA20,0x%h_0x%h\n0xEA40,0x%h_0x%h\n0xEA60,0x%h_0x%h\n0xEA80,0x%h_0x%h\n0xEAA0,0x%h_0x%h\n0xEAC0,0x%h_0x%h\n0xEAE0,0x%h_0x%h\n0xEB00,0x%h_0x%h\n0xEB20,0x%h_0x%h\n0xEB40,0x%h_0x%h\n0xEB60,0x%h_0x%h\n0xEB80,0x%h_0x%h\n0xEBA0,0x%h_0x%h\n0xEBC0,0x%h_0x%h\n0xEBE0,0x%h_0x%h\n0xEC00,0x%h_0x%h\n0xEC20,0x%h_0x%h\n0xEC40,0x%h_0x%h\n0xEC60,0x%h_0x%h\n0xEC80,0x%h_0x%h\n0xECA0,0x%h_0x%h\n0xECC0,0x%h_0x%h\n0xECE0,0x%h_0x%h\n0xED00,0x%h_0x%h\n0xED20,0x%h_0x%h\n0xED40,0x%h_0x%h\n0xED60,0x%h_0x%h\n0xED80,0x%h_0x%h\n0xEDA0,0x%h_0x%h\n0xEDC0,0x%h_0x%h\n0xEDE0,0x%h_0x%h\n0xEE00,0x%h_0x%h\n0xEE20,0x%h_0x%h\n0xEE40,0x%h_0x%h\n0xEE60,0x%h_0x%h\n0xEE80,0x%h_0x%h\n0xEEA0,0x%h_0x%h\n0xEEC0,0x%h_0x%h\n0xEEE0,0x%h_0x%h\n0xEF00,0x%h_0x%h\n0xEF20,0x%h_0x%h\n0xEF40,0x%h_0x%h\n0xEF60,0x%h_0x%h\n0xEF80,0x%h_0x%h\n0xEFA0,0x%h_0x%h\n0xEFC0,0x%h_0x%h\n0xEFE0,0x%h_0x%h\n0xF000,0x%h_0x%h\n0xF020,0x%h_0x%h\n0xF040,0x%h_0x%h\n0xF060,0x%h_0x%h\n0xF080,0x%h_0x%h\n0xF0A0,0x%h_0x%h\n0xF0C0,0x%h_0x%h\n0xF0E0,0x%h_0x%h\n0xF100,0x%h_0x%h\n0xF120,0x%h_0x%h\n0xF140,0x%h_0x%h\n0xF160,0x%h_0x%h\n0xF180,0x%h_0x%h\n0xF1A0,0x%h_0x%h\n0xF1C0,0x%h_0x%h\n0xF1E0,0x%h_0x%h\n0xF200,0x%h_0x%h\n0xF220,0x%h_0x%h\n0xF240,0x%h_0x%h\n0xF260,0x%h_0x%h\n0xF280,0x%h_0x%h\n0xF2A0,0x%h_0x%h\n0xF2C0,0x%h_0x%h\n0xF2E0,0x%h_0x%h\n0xF300,0x%h_0x%h\n0xF320,0x%h_0x%h\n0xF340,0x%h_0x%h\n0xF360,0x%h_0x%h\n0xF380,0x%h_0x%h\n0xF3A0,0x%h_0x%h\n0xF3C0,0x%h_0x%h\n0xF3E0,0x%h_0x%h\n0xF400,0x%h_0x%h\n0xF420,0x%h_0x%h\n0xF440,0x%h_0x%h\n0xF460,0x%h_0x%h\n0xF480,0x%h_0x%h\n0xF4A0,0x%h_0x%h\n0xF4C0,0x%h_0x%h\n0xF4E0,0x%h_0x%h\n0xF500,0x%h_0x%h\n0xF520,0x%h_0x%h\n0xF540,0x%h_0x%h\n0xF560,0x%h_0x%h\n0xF580,0x%h_0x%h\n0xF5A0,0x%h_0x%h\n0xF5C0,0x%h_0x%h\n0xF5E0,0x%h_0x%h\n0xF600,0x%h_0x%h\n0xF620,0x%h_0x%h\n0xF640,0x%h_0x%h\n0xF660,0x%h_0x%h\n0xF680,0x%h_0x%h\n0xF6A0,0x%h_0x%h\n0xF6C0,0x%h_0x%h\n0xF6E0,0x%h_0x%h\n0xF700,0x%h_0x%h\n0xF720,0x%h_0x%h\n0xF740,0x%h_0x%h\n0xF760,0x%h_0x%h\n0xF780,0x%h_0x%h\n0xF7A0,0x%h_0x%h\n0xF7C0,0x%h_0x%h\n0xF7E0,0x%h_0x%h\n0xF800,0x%h_0x%h\n0xF820,0x%h_0x%h\n0xF840,0x%h_0x%h\n0xF860,0x%h_0x%h\n0xF880,0x%h_0x%h\n0xF8A0,0x%h_0x%h\n0xF8C0,0x%h_0x%h\n0xF8E0,0x%h_0x%h\n0xF900,0x%h_0x%h\n0xF920,0x%h_0x%h\n0xF940,0x%h_0x%h\n0xF960,0x%h_0x%h\n0xF980,0x%h_0x%h\n0xF9A0,0x%h_0x%h\n0xF9C0,0x%h_0x%h\n0xF9E0,0x%h_0x%h\n0xFA00,0x%h_0x%h\n0xFA20,0x%h_0x%h\n0xFA40,0x%h_0x%h\n0xFA60,0x%h_0x%h\n0xFA80,0x%h_0x%h\n0xFAA0,0x%h_0x%h\n0xFAC0,0x%h_0x%h\n0xFAE0,0x%h_0x%h\n0xFB00,0x%h_0x%h\n0xFB20,0x%h_0x%h\n0xFB40,0x%h_0x%h\n0xFB60,0x%h_0x%h\n0xFB80,0x%h_0x%h\n0xFBA0,0x%h_0x%h\n0xFBC0,0x%h_0x%h\n0xFBE0,0x%h_0x%h\n0xFC00,0x%h_0x%h\n0xFC20,0x%h_0x%h\n0xFC40,0x%h_0x%h\n0xFC60,0x%h_0x%h\n0xFC80,0x%h_0x%h\n0xFCA0,0x%h_0x%h\n0xFCC0,0x%h_0x%h\n0xFCE0,0x%h_0x%h\n0xFD00,0x%h_0x%h\n0xFD20,0x%h_0x%h\n0xFD40,0x%h_0x%h\n0xFD60,0x%h_0x%h\n0xFD80,0x%h_0x%h\n0xFDA0,0x%h_0x%h\n0xFDC0,0x%h_0x%h\n0xFDE0,0x%h_0x%h\n0xFE00,0x%h_0x%h\n0xFE20,0x%h_0x%h\n0xFE40,0x%h_0x%h\n0xFE60,0x%h_0x%h\n0xFE80,0x%h_0x%h\n0xFEA0,0x%h_0x%h\n0xFEC0,0x%h_0x%h\n0xFEE0,0x%h_0x%h\n0xFF00,0x%h_0x%h\n0xFF20,0x%h_0x%h\n0xFF40,0x%h_0x%h\n0xFF60,0x%h_0x%h\n0xFF80,0x%h_0x%h\n0xFFA0,0x%h_0x%h\n0xFFC0,0x%h_0x%h\n0xFFE0,0x%h_0x%h\n0x10000,0x%h_0x%h\n0x10020,0x%h_0x%h\n0x10040,0x%h_0x%h\n0x10060,0x%h_0x%h\n0x10080,0x%h_0x%h\n0x100A0,0x%h_0x%h\n0x100C0,0x%h_0x%h\n0x100E0,0x%h_0x%h\n0x10100,0x%h_0x%h\n0x10120,0x%h_0x%h\n0x10140,0x%h_0x%h\n0x10160,0x%h_0x%h\n0x10180,0x%h_0x%h\n0x101A0,0x%h_0x%h\n0x101C0,0x%h_0x%h\n0x101E0,0x%h_0x%h\n0x10200,0x%h_0x%h\n0x10220,0x%h_0x%h\n0x10240,0x%h_0x%h\n0x10260,0x%h_0x%h\n0x10280,0x%h_0x%h\n0x102A0,0x%h_0x%h\n0x102C0,0x%h_0x%h\n0x102E0,0x%h_0x%h\n0x10300,0x%h_0x%h\n0x10320,0x%h_0x%h\n0x10340,0x%h_0x%h\n0x10360,0x%h_0x%h\n0x10380,0x%h_0x%h\n0x103A0,0x%h_0x%h\n0x103C0,0x%h_0x%h\n0x103E0,0x%h_0x%h\n0x10400,0x%h_0x%h\n0x10420,0x%h_0x%h\n0x10440,0x%h_0x%h\n0x10460,0x%h_0x%h\n0x10480,0x%h_0x%h\n0x104A0,0x%h_0x%h\n0x104C0,0x%h_0x%h\n0x104E0,0x%h_0x%h\n0x10500,0x%h_0x%h\n0x10520,0x%h_0x%h\n0x10540,0x%h_0x%h\n0x10560,0x%h_0x%h\n0x10580,0x%h_0x%h\n0x105A0,0x%h_0x%h\n0x105C0,0x%h_0x%h\n0x105E0,0x%h_0x%h\n0x10600,0x%h_0x%h\n0x10620,0x%h_0x%h\n0x10640,0x%h_0x%h\n0x10660,0x%h_0x%h\n0x10680,0x%h_0x%h\n0x106A0,0x%h_0x%h\n0x106C0,0x%h_0x%h\n0x106E0,0x%h_0x%h\n0x10700,0x%h_0x%h\n0x10720,0x%h_0x%h\n0x10740,0x%h_0x%h\n0x10760,0x%h_0x%h\n0x10780,0x%h_0x%h\n0x107A0,0x%h_0x%h\n0x107C0,0x%h_0x%h\n0x107E0,0x%h_0x%h\n0x10800,0x%h_0x%h\n0x10820,0x%h_0x%h\n0x10840,0x%h_0x%h\n0x10860,0x%h_0x%h\n0x10880,0x%h_0x%h\n0x108A0,0x%h_0x%h\n0x108C0,0x%h_0x%h\n0x108E0,0x%h_0x%h\n0x10900,0x%h_0x%h\n0x10920,0x%h_0x%h\n0x10940,0x%h_0x%h\n0x10960,0x%h_0x%h\n0x10980,0x%h_0x%h\n0x109A0,0x%h_0x%h\n0x109C0,0x%h_0x%h\n0x109E0,0x%h_0x%h\n0x10A00,0x%h_0x%h\n0x10A20,0x%h_0x%h\n0x10A40,0x%h_0x%h\n0x10A60,0x%h_0x%h\n0x10A80,0x%h_0x%h\n0x10AA0,0x%h_0x%h\n0x10AC0,0x%h_0x%h\n0x10AE0,0x%h_0x%h\n0x10B00,0x%h_0x%h\n0x10B20,0x%h_0x%h\n0x10B40,0x%h_0x%h\n0x10B60,0x%h_0x%h\n0x10B80,0x%h_0x%h\n0x10BA0,0x%h_0x%h\n0x10BC0,0x%h_0x%h\n0x10BE0,0x%h_0x%h\n0x10C00,0x%h_0x%h\n0x10C20,0x%h_0x%h\n0x10C40,0x%h_0x%h\n0x10C60,0x%h_0x%h\n0x10C80,0x%h_0x%h\n0x10CA0,0x%h_0x%h\n0x10CC0,0x%h_0x%h\n0x10CE0,0x%h_0x%h\n0x10D00,0x%h_0x%h\n0x10D20,0x%h_0x%h\n0x10D40,0x%h_0x%h\n0x10D60,0x%h_0x%h\n0x10D80,0x%h_0x%h\n0x10DA0,0x%h_0x%h\n0x10DC0,0x%h_0x%h\n0x10DE0,0x%h_0x%h\n0x10E00,0x%h_0x%h\n0x10E20,0x%h_0x%h\n0x10E40,0x%h_0x%h\n0x10E60,0x%h_0x%h\n0x10E80,0x%h_0x%h\n0x10EA0,0x%h_0x%h\n0x10EC0,0x%h_0x%h\n0x10EE0,0x%h_0x%h\n0x10F00,0x%h_0x%h\n0x10F20,0x%h_0x%h\n0x10F40,0x%h_0x%h\n0x10F60,0x%h_0x%h\n0x10F80,0x%h_0x%h\n0x10FA0,0x%h_0x%h\n0x10FC0,0x%h_0x%h\n0x10FE0,0x%h_0x%h\n0x11000,0x%h_0x%h\n0x11020,0x%h_0x%h\n0x11040,0x%h_0x%h\n0x11060,0x%h_0x%h\n0x11080,0x%h_0x%h\n0x110A0,0x%h_0x%h\n0x110C0,0x%h_0x%h\n0x110E0,0x%h_0x%h\n0x11100,0x%h_0x%h\n0x11120,0x%h_0x%h\n0x11140,0x%h_0x%h\n0x11160,0x%h_0x%h\n0x11180,0x%h_0x%h\n0x111A0,0x%h_0x%h\n0x111C0,0x%h_0x%h\n0x111E0,0x%h_0x%h\n0x11200,0x%h_0x%h\n0x11220,0x%h_0x%h\n0x11240,0x%h_0x%h\n0x11260,0x%h_0x%h\n0x11280,0x%h_0x%h\n0x112A0,0x%h_0x%h\n0x112C0,0x%h_0x%h\n0x112E0,0x%h_0x%h\n0x11300,0x%h_0x%h\n0x11320,0x%h_0x%h\n0x11340,0x%h_0x%h\n0x11360,0x%h_0x%h\n0x11380,0x%h_0x%h\n0x113A0,0x%h_0x%h\n0x113C0,0x%h_0x%h\n0x113E0,0x%h_0x%h\n0x11400,0x%h_0x%h\n0x11420,0x%h_0x%h\n0x11440,0x%h_0x%h\n0x11460,0x%h_0x%h\n0x11480,0x%h_0x%h\n0x114A0,0x%h_0x%h\n0x114C0,0x%h_0x%h\n0x114E0,0x%h_0x%h\n0x11500,0x%h_0x%h\n0x11520,0x%h_0x%h\n0x11540,0x%h_0x%h\n0x11560,0x%h_0x%h\n0x11580,0x%h_0x%h\n0x115A0,0x%h_0x%h\n0x115C0,0x%h_0x%h\n0x115E0,0x%h_0x%h\n0x11600,0x%h_0x%h\n0x11620,0x%h_0x%h\n0x11640,0x%h_0x%h\n0x11660,0x%h_0x%h\n0x11680,0x%h_0x%h\n0x116A0,0x%h_0x%h\n0x116C0,0x%h_0x%h\n0x116E0,0x%h_0x%h\n0x11700,0x%h_0x%h\n0x11720,0x%h_0x%h\n0x11740,0x%h_0x%h\n0x11760,0x%h_0x%h\n0x11780,0x%h_0x%h\n0x117A0,0x%h_0x%h\n0x117C0,0x%h_0x%h\n0x117E0,0x%h_0x%h\n0x11800,0x%h_0x%h\n0x11820,0x%h_0x%h\n0x11840,0x%h_0x%h\n0x11860,0x%h_0x%h\n0x11880,0x%h_0x%h\n0x118A0,0x%h_0x%h\n0x118C0,0x%h_0x%h\n0x118E0,0x%h_0x%h\n0x11900,0x%h_0x%h\n0x11920,0x%h_0x%h\n0x11940,0x%h_0x%h\n0x11960,0x%h_0x%h\n0x11980,0x%h_0x%h\n0x119A0,0x%h_0x%h\n0x119C0,0x%h_0x%h\n0x119E0,0x%h_0x%h\n0x11A00,0x%h_0x%h\n0x11A20,0x%h_0x%h\n0x11A40,0x%h_0x%h\n0x11A60,0x%h_0x%h\n0x11A80,0x%h_0x%h\n0x11AA0,0x%h_0x%h\n0x11AC0,0x%h_0x%h\n0x11AE0,0x%h_0x%h\n0x11B00,0x%h_0x%h\n0x11B20,0x%h_0x%h\n0x11B40,0x%h_0x%h\n0x11B60,0x%h_0x%h\n0x11B80,0x%h_0x%h\n0x11BA0,0x%h_0x%h\n0x11BC0,0x%h_0x%h\n0x11BE0,0x%h_0x%h\n0x11C00,0x%h_0x%h\n0x11C20,0x%h_0x%h\n0x11C40,0x%h_0x%h\n0x11C60,0x%h_0x%h\n0x11C80,0x%h_0x%h\n0x11CA0,0x%h_0x%h\n0x11CC0,0x%h_0x%h\n0x11CE0,0x%h_0x%h\n0x11D00,0x%h_0x%h\n0x11D20,0x%h_0x%h\n0x11D40,0x%h_0x%h\n0x11D60,0x%h_0x%h\n0x11D80,0x%h_0x%h\n0x11DA0,0x%h_0x%h\n0x11DC0,0x%h_0x%h\n0x11DE0,0x%h_0x%h\n0x11E00,0x%h_0x%h\n0x11E20,0x%h_0x%h\n0x11E40,0x%h_0x%h\n0x11E60,0x%h_0x%h\n0x11E80,0x%h_0x%h\n0x11EA0,0x%h_0x%h\n0x11EC0,0x%h_0x%h\n0x11EE0,0x%h_0x%h\n0x11F00,0x%h_0x%h\n0x11F20,0x%h_0x%h\n0x11F40,0x%h_0x%h\n0x11F60,0x%h_0x%h\n0x11F80,0x%h_0x%h\n0x11FA0,0x%h_0x%h\n0x11FC0,0x%h_0x%h\n0x11FE0,0x%h_0x%h\n0x12000,0x%h_0x%h\n0x12020,0x%h_0x%h\n0x12040,0x%h_0x%h\n0x12060,0x%h_0x%h\n0x12080,0x%h_0x%h\n0x120A0,0x%h_0x%h\n0x120C0,0x%h_0x%h\n0x120E0,0x%h_0x%h\n0x12100,0x%h_0x%h\n0x12120,0x%h_0x%h\n0x12140,0x%h_0x%h\n0x12160,0x%h_0x%h\n0x12180,0x%h_0x%h\n0x121A0,0x%h_0x%h\n0x121C0,0x%h_0x%h\n0x121E0,0x%h_0x%h\n0x12200,0x%h_0x%h\n0x12220,0x%h_0x%h\n0x12240,0x%h_0x%h\n0x12260,0x%h_0x%h\n0x12280,0x%h_0x%h\n0x122A0,0x%h_0x%h\n0x122C0,0x%h_0x%h\n0x122E0,0x%h_0x%h\n0x12300,0x%h_0x%h\n0x12320,0x%h_0x%h\n0x12340,0x%h_0x%h\n0x12360,0x%h_0x%h\n0x12380,0x%h_0x%h\n0x123A0,0x%h_0x%h\n0x123C0,0x%h_0x%h\n0x123E0,0x%h_0x%h\n0x12400,0x%h_0x%h\n0x12420,0x%h_0x%h\n0x12440,0x%h_0x%h\n0x12460,0x%h_0x%h\n0x12480,0x%h_0x%h\n0x124A0,0x%h_0x%h\n0x124C0,0x%h_0x%h\n0x124E0,0x%h_0x%h\n0x12500,0x%h_0x%h\n0x12520,0x%h_0x%h\n0x12540,0x%h_0x%h\n0x12560,0x%h_0x%h\n0x12580,0x%h_0x%h\n0x125A0,0x%h_0x%h\n0x125C0,0x%h_0x%h\n0x125E0,0x%h_0x%h\n0x12600,0x%h_0x%h\n0x12620,0x%h_0x%h\n0x12640,0x%h_0x%h\n0x12660,0x%h_0x%h\n0x12680,0x%h_0x%h\n0x126A0,0x%h_0x%h\n0x126C0,0x%h_0x%h\n0x126E0,0x%h_0x%h\n0x12700,0x%h_0x%h\n0x12720,0x%h_0x%h\n0x12740,0x%h_0x%h\n0x12760,0x%h_0x%h\n0x12780,0x%h_0x%h\n0x127A0,0x%h_0x%h\n0x127C0,0x%h_0x%h\n0x127E0,0x%h_0x%h\n0x12800,0x%h_0x%h\n0x12820,0x%h_0x%h\n0x12840,0x%h_0x%h\n0x12860,0x%h_0x%h\n0x12880,0x%h_0x%h\n0x128A0,0x%h_0x%h\n0x128C0,0x%h_0x%h\n0x128E0,0x%h_0x%h\n0x12900,0x%h_0x%h\n0x12920,0x%h_0x%h\n0x12940,0x%h_0x%h\n0x12960,0x%h_0x%h\n0x12980,0x%h_0x%h\n0x129A0,0x%h_0x%h\n0x129C0,0x%h_0x%h\n0x129E0,0x%h_0x%h\n0x12A00,0x%h_0x%h\n0x12A20,0x%h_0x%h\n0x12A40,0x%h_0x%h\n0x12A60,0x%h_0x%h\n0x12A80,0x%h_0x%h\n0x12AA0,0x%h_0x%h\n0x12AC0,0x%h_0x%h\n0x12AE0,0x%h_0x%h\n0x12B00,0x%h_0x%h\n0x12B20,0x%h_0x%h\n0x12B40,0x%h_0x%h\n0x12B60,0x%h_0x%h\n0x12B80,0x%h_0x%h\n0x12BA0,0x%h_0x%h\n0x12BC0,0x%h_0x%h\n0x12BE0,0x%h_0x%h\n0x12C00,0x%h_0x%h\n0x12C20,0x%h_0x%h\n0x12C40,0x%h_0x%h\n0x12C60,0x%h_0x%h\n0x12C80,0x%h_0x%h\n0x12CA0,0x%h_0x%h\n0x12CC0,0x%h_0x%h\n0x12CE0,0x%h_0x%h\n0x12D00,0x%h_0x%h\n0x12D20,0x%h_0x%h\n0x12D40,0x%h_0x%h\n0x12D60,0x%h_0x%h\n0x12D80,0x%h_0x%h\n0x12DA0,0x%h_0x%h\n0x12DC0,0x%h_0x%h\n0x12DE0,0x%h_0x%h\n0x12E00,0x%h_0x%h\n0x12E20,0x%h_0x%h\n0x12E40,0x%h_0x%h\n0x12E60,0x%h_0x%h\n0x12E80,0x%h_0x%h\n0x12EA0,0x%h_0x%h\n0x12EC0,0x%h_0x%h\n0x12EE0,0x%h_0x%h\n0x12F00,0x%h_0x%h\n0x12F20,0x%h_0x%h\n0x12F40,0x%h_0x%h\n0x12F60,0x%h_0x%h\n0x12F80,0x%h_0x%h\n0x12FA0,0x%h_0x%h\n0x12FC0,0x%h_0x%h\n0x12FE0,0x%h_0x%h\n0x13000,0x%h_0x%h\n0x13020,0x%h_0x%h\n0x13040,0x%h_0x%h\n0x13060,0x%h_0x%h\n0x13080,0x%h_0x%h\n0x130A0,0x%h_0x%h\n0x130C0,0x%h_0x%h\n0x130E0,0x%h_0x%h\n0x13100,0x%h_0x%h\n0x13120,0x%h_0x%h\n0x13140,0x%h_0x%h\n0x13160,0x%h_0x%h\n0x13180,0x%h_0x%h\n0x131A0,0x%h_0x%h\n0x131C0,0x%h_0x%h\n0x131E0,0x%h_0x%h\n0x13200,0x%h_0x%h\n0x13220,0x%h_0x%h\n0x13240,0x%h_0x%h\n0x13260,0x%h_0x%h\n0x13280,0x%h_0x%h\n0x132A0,0x%h_0x%h\n0x132C0,0x%h_0x%h\n0x132E0,0x%h_0x%h\n0x13300,0x%h_0x%h\n0x13320,0x%h_0x%h\n0x13340,0x%h_0x%h\n0x13360,0x%h_0x%h\n0x13380,0x%h_0x%h\n0x133A0,0x%h_0x%h\n0x133C0,0x%h_0x%h\n0x133E0,0x%h_0x%h\n0x13400,0x%h_0x%h\n0x13420,0x%h_0x%h\n0x13440,0x%h_0x%h\n0x13460,0x%h_0x%h\n0x13480,0x%h_0x%h\n0x134A0,0x%h_0x%h\n0x134C0,0x%h_0x%h\n0x134E0,0x%h_0x%h\n0x13500,0x%h_0x%h\n0x13520,0x%h_0x%h\n0x13540,0x%h_0x%h\n0x13560,0x%h_0x%h\n0x13580,0x%h_0x%h\n0x135A0,0x%h_0x%h\n0x135C0,0x%h_0x%h\n0x135E0,0x%h_0x%h\n0x13600,0x%h_0x%h\n0x13620,0x%h_0x%h\n0x13640,0x%h_0x%h\n0x13660,0x%h_0x%h\n0x13680,0x%h_0x%h\n0x136A0,0x%h_0x%h\n0x136C0,0x%h_0x%h\n0x136E0,0x%h_0x%h\n0x13700,0x%h_0x%h\n0x13720,0x%h_0x%h\n0x13740,0x%h_0x%h\n0x13760,0x%h_0x%h\n0x13780,0x%h_0x%h\n0x137A0,0x%h_0x%h\n0x137C0,0x%h_0x%h\n0x137E0,0x%h_0x%h\n0x13800,0x%h_0x%h\n0x13820,0x%h_0x%h\n0x13840,0x%h_0x%h\n0x13860,0x%h_0x%h\n0x13880,0x%h_0x%h\n0x138A0,0x%h_0x%h\n0x138C0,0x%h_0x%h\n0x138E0,0x%h_0x%h\n0x13900,0x%h_0x%h\n0x13920,0x%h_0x%h\n0x13940,0x%h_0x%h\n0x13960,0x%h_0x%h\n0x13980,0x%h_0x%h\n0x139A0,0x%h_0x%h\n0x139C0,0x%h_0x%h\n0x139E0,0x%h_0x%h\n0x13A00,0x%h_0x%h\n0x13A20,0x%h_0x%h\n0x13A40,0x%h_0x%h\n0x13A60,0x%h_0x%h\n0x13A80,0x%h_0x%h\n0x13AA0,0x%h_0x%h\n0x13AC0,0x%h_0x%h\n0x13AE0,0x%h_0x%h\n0x13B00,0x%h_0x%h\n0x13B20,0x%h_0x%h\n0x13B40,0x%h_0x%h\n0x13B60,0x%h_0x%h\n0x13B80,0x%h_0x%h\n0x13BA0,0x%h_0x%h\n0x13BC0,0x%h_0x%h\n0x13BE0,0x%h_0x%h\n0x13C00,0x%h_0x%h\n0x13C20,0x%h_0x%h\n0x13C40,0x%h_0x%h\n0x13C60,0x%h_0x%h\n0x13C80,0x%h_0x%h\n0x13CA0,0x%h_0x%h\n0x13CC0,0x%h_0x%h\n0x13CE0,0x%h_0x%h\n0x13D00,0x%h_0x%h\n0x13D20,0x%h_0x%h\n0x13D40,0x%h_0x%h\n0x13D60,0x%h_0x%h\n0x13D80,0x%h_0x%h\n0x13DA0,0x%h_0x%h\n0x13DC0,0x%h_0x%h\n0x13DE0,0x%h_0x%h\n0x13E00,0x%h_0x%h\n0x13E20,0x%h_0x%h\n0x13E40,0x%h_0x%h\n0x13E60,0x%h_0x%h\n0x13E80,0x%h_0x%h\n0x13EA0,0x%h_0x%h\n0x13EC0,0x%h_0x%h\n0x13EE0,0x%h_0x%h\n0x13F00,0x%h_0x%h\n0x13F20,0x%h_0x%h\n0x13F40,0x%h_0x%h\n0x13F60,0x%h_0x%h\n0x13F80,0x%h_0x%h\n0x13FA0,0x%h_0x%h\n0x13FC0,0x%h_0x%h\n0x13FE0,0x%h_0x%h\n0x14000,0x%h_0x%h\n0x14020,0x%h_0x%h\n0x14040,0x%h_0x%h\n0x14060,0x%h_0x%h\n0x14080,0x%h_0x%h\n0x140A0,0x%h_0x%h\n0x140C0,0x%h_0x%h\n0x140E0,0x%h_0x%h\n0x14100,0x%h_0x%h\n0x14120,0x%h_0x%h\n0x14140,0x%h_0x%h\n0x14160,0x%h_0x%h\n0x14180,0x%h_0x%h\n0x141A0,0x%h_0x%h\n0x141C0,0x%h_0x%h\n0x141E0,0x%h_0x%h\n0x14200,0x%h_0x%h\n0x14220,0x%h_0x%h\n0x14240,0x%h_0x%h\n0x14260,0x%h_0x%h\n0x14280,0x%h_0x%h\n0x142A0,0x%h_0x%h\n0x142C0,0x%h_0x%h\n0x142E0,0x%h_0x%h\n0x14300,0x%h_0x%h\n0x14320,0x%h_0x%h\n0x14340,0x%h_0x%h\n0x14360,0x%h_0x%h\n0x14380,0x%h_0x%h\n0x143A0,0x%h_0x%h\n0x143C0,0x%h_0x%h\n0x143E0,0x%h_0x%h\n0x14400,0x%h_0x%h\n0x14420,0x%h_0x%h\n0x14440,0x%h_0x%h\n0x14460,0x%h_0x%h\n0x14480,0x%h_0x%h\n0x144A0,0x%h_0x%h\n0x144C0,0x%h_0x%h\n0x144E0,0x%h_0x%h\n0x14500,0x%h_0x%h\n0x14520,0x%h_0x%h\n0x14540,0x%h_0x%h\n0x14560,0x%h_0x%h\n0x14580,0x%h_0x%h\n0x145A0,0x%h_0x%h\n0x145C0,0x%h_0x%h\n0x145E0,0x%h_0x%h\n0x14600,0x%h_0x%h\n0x14620,0x%h_0x%h\n0x14640,0x%h_0x%h\n0x14660,0x%h_0x%h\n0x14680,0x%h_0x%h\n0x146A0,0x%h_0x%h\n0x146C0,0x%h_0x%h\n0x146E0,0x%h_0x%h\n0x14700,0x%h_0x%h\n0x14720,0x%h_0x%h\n0x14740,0x%h_0x%h\n0x14760,0x%h_0x%h\n0x14780,0x%h_0x%h\n0x147A0,0x%h_0x%h\n0x147C0,0x%h_0x%h\n0x147E0,0x%h_0x%h\n0x14800,0x%h_0x%h\n0x14820,0x%h_0x%h\n0x14840,0x%h_0x%h\n0x14860,0x%h_0x%h\n0x14880,0x%h_0x%h\n0x148A0,0x%h_0x%h\n0x148C0,0x%h_0x%h\n0x148E0,0x%h_0x%h\n0x14900,0x%h_0x%h\n0x14920,0x%h_0x%h\n0x14940,0x%h_0x%h\n0x14960,0x%h_0x%h\n0x14980,0x%h_0x%h\n0x149A0,0x%h_0x%h\n0x149C0,0x%h_0x%h\n0x149E0,0x%h_0x%h\n0x14A00,0x%h_0x%h\n0x14A20,0x%h_0x%h\n0x14A40,0x%h_0x%h\n0x14A60,0x%h_0x%h\n0x14A80,0x%h_0x%h\n0x14AA0,0x%h_0x%h\n0x14AC0,0x%h_0x%h\n0x14AE0,0x%h_0x%h\n0x14B00,0x%h_0x%h\n0x14B20,0x%h_0x%h\n0x14B40,0x%h_0x%h\n0x14B60,0x%h_0x%h\n0x14B80,0x%h_0x%h\n0x14BA0,0x%h_0x%h\n0x14BC0,0x%h_0x%h\n0x14BE0,0x%h_0x%h\n0x14C00,0x%h_0x%h\n0x14C20,0x%h_0x%h\n0x14C40,0x%h_0x%h\n0x14C60,0x%h_0x%h\n0x14C80,0x%h_0x%h\n0x14CA0,0x%h_0x%h\n0x14CC0,0x%h_0x%h\n0x14CE0,0x%h_0x%h\n0x14D00,0x%h_0x%h\n0x14D20,0x%h_0x%h\n0x14D40,0x%h_0x%h\n0x14D60,0x%h_0x%h\n0x14D80,0x%h_0x%h\n0x14DA0,0x%h_0x%h\n0x14DC0,0x%h_0x%h\n0x14DE0,0x%h_0x%h\n0x14E00,0x%h_0x%h\n0x14E20,0x%h_0x%h\n0x14E40,0x%h_0x%h\n0x14E60,0x%h_0x%h\n0x14E80,0x%h_0x%h\n0x14EA0,0x%h_0x%h\n0x14EC0,0x%h_0x%h\n0x14EE0,0x%h_0x%h\n0x14F00,0x%h_0x%h\n0x14F20,0x%h_0x%h\n0x14F40,0x%h_0x%h\n0x14F60,0x%h_0x%h\n0x14F80,0x%h_0x%h\n0x14FA0,0x%h_0x%h\n0x14FC0,0x%h_0x%h\n0x14FE0,0x%h_0x%h\n0x15000,0x%h_0x%h\n0x15020,0x%h_0x%h\n0x15040,0x%h_0x%h\n0x15060,0x%h_0x%h\n0x15080,0x%h_0x%h\n0x150A0,0x%h_0x%h\n0x150C0,0x%h_0x%h\n0x150E0,0x%h_0x%h\n0x15100,0x%h_0x%h\n0x15120,0x%h_0x%h\n0x15140,0x%h_0x%h\n0x15160,0x%h_0x%h\n0x15180,0x%h_0x%h\n0x151A0,0x%h_0x%h\n0x151C0,0x%h_0x%h\n0x151E0,0x%h_0x%h\n0x15200,0x%h_0x%h\n0x15220,0x%h_0x%h\n0x15240,0x%h_0x%h\n0x15260,0x%h_0x%h\n0x15280,0x%h_0x%h\n0x152A0,0x%h_0x%h\n0x152C0,0x%h_0x%h\n0x152E0,0x%h_0x%h\n0x15300,0x%h_0x%h\n0x15320,0x%h_0x%h\n0x15340,0x%h_0x%h\n0x15360,0x%h_0x%h\n0x15380,0x%h_0x%h\n0x153A0,0x%h_0x%h\n0x153C0,0x%h_0x%h\n0x153E0,0x%h_0x%h\n0x15400,0x%h_0x%h\n0x15420,0x%h_0x%h\n0x15440,0x%h_0x%h\n0x15460,0x%h_0x%h\n0x15480,0x%h_0x%h\n0x154A0,0x%h_0x%h\n0x154C0,0x%h_0x%h\n0x154E0,0x%h_0x%h\n0x15500,0x%h_0x%h\n0x15520,0x%h_0x%h\n0x15540,0x%h_0x%h\n0x15560,0x%h_0x%h\n0x15580,0x%h_0x%h\n0x155A0,0x%h_0x%h\n0x155C0,0x%h_0x%h\n0x155E0,0x%h_0x%h\n0x15600,0x%h_0x%h\n0x15620,0x%h_0x%h\n0x15640,0x%h_0x%h\n0x15660,0x%h_0x%h\n0x15680,0x%h_0x%h\n0x156A0,0x%h_0x%h\n0x156C0,0x%h_0x%h\n0x156E0,0x%h_0x%h\n0x15700,0x%h_0x%h\n0x15720,0x%h_0x%h\n0x15740,0x%h_0x%h\n0x15760,0x%h_0x%h\n0x15780,0x%h_0x%h\n0x157A0,0x%h_0x%h\n0x157C0,0x%h_0x%h\n0x157E0,0x%h_0x%h\n0x15800,0x%h_0x%h\n0x15820,0x%h_0x%h\n0x15840,0x%h_0x%h\n0x15860,0x%h_0x%h\n0x15880,0x%h_0x%h\n0x158A0,0x%h_0x%h\n0x158C0,0x%h_0x%h\n0x158E0,0x%h_0x%h\n0x15900,0x%h_0x%h\n0x15920,0x%h_0x%h\n0x15940,0x%h_0x%h\n0x15960,0x%h_0x%h\n0x15980,0x%h_0x%h\n0x159A0,0x%h_0x%h\n0x159C0,0x%h_0x%h\n0x159E0,0x%h_0x%h\n0x15A00,0x%h_0x%h\n0x15A20,0x%h_0x%h\n0x15A40,0x%h_0x%h\n0x15A60,0x%h_0x%h\n0x15A80,0x%h_0x%h\n0x15AA0,0x%h_0x%h\n0x15AC0,0x%h_0x%h\n0x15AE0,0x%h_0x%h\n0x15B00,0x%h_0x%h\n0x15B20,0x%h_0x%h\n0x15B40,0x%h_0x%h\n0x15B60,0x%h_0x%h\n0x15B80,0x%h_0x%h\n0x15BA0,0x%h_0x%h\n0x15BC0,0x%h_0x%h\n0x15BE0,0x%h_0x%h\n0x15C00,0x%h_0x%h\n0x15C20,0x%h_0x%h\n0x15C40,0x%h_0x%h\n0x15C60,0x%h_0x%h\n0x15C80,0x%h_0x%h\n0x15CA0,0x%h_0x%h\n0x15CC0,0x%h_0x%h\n0x15CE0,0x%h_0x%h\n0x15D00,0x%h_0x%h\n0x15D20,0x%h_0x%h\n0x15D40,0x%h_0x%h\n0x15D60,0x%h_0x%h\n0x15D80,0x%h_0x%h\n0x15DA0,0x%h_0x%h\n0x15DC0,0x%h_0x%h\n0x15DE0,0x%h_0x%h\n0x15E00,0x%h_0x%h\n0x15E20,0x%h_0x%h\n0x15E40,0x%h_0x%h\n0x15E60,0x%h_0x%h\n0x15E80,0x%h_0x%h\n0x15EA0,0x%h_0x%h\n0x15EC0,0x%h_0x%h\n0x15EE0,0x%h_0x%h\n0x15F00,0x%h_0x%h\n0x15F20,0x%h_0x%h\n0x15F40,0x%h_0x%h\n0x15F60,0x%h_0x%h\n0x15F80,0x%h_0x%h\n0x15FA0,0x%h_0x%h\n0x15FC0,0x%h_0x%h\n0x15FE0,0x%h_0x%h\n0x16000,0x%h_0x%h\n0x16020,0x%h_0x%h\n0x16040,0x%h_0x%h\n0x16060,0x%h_0x%h\n0x16080,0x%h_0x%h\n0x160A0,0x%h_0x%h\n0x160C0,0x%h_0x%h\n0x160E0,0x%h_0x%h\n0x16100,0x%h_0x%h\n0x16120,0x%h_0x%h\n0x16140,0x%h_0x%h\n0x16160,0x%h_0x%h\n0x16180,0x%h_0x%h\n0x161A0,0x%h_0x%h\n0x161C0,0x%h_0x%h\n0x161E0,0x%h_0x%h\n0x16200,0x%h_0x%h\n0x16220,0x%h_0x%h\n0x16240,0x%h_0x%h\n0x16260,0x%h_0x%h\n0x16280,0x%h_0x%h\n0x162A0,0x%h_0x%h\n0x162C0,0x%h_0x%h\n0x162E0,0x%h_0x%h\n0x16300,0x%h_0x%h\n0x16320,0x%h_0x%h\n0x16340,0x%h_0x%h\n0x16360,0x%h_0x%h\n0x16380,0x%h_0x%h\n0x163A0,0x%h_0x%h\n0x163C0,0x%h_0x%h\n0x163E0,0x%h_0x%h\n0x16400,0x%h_0x%h\n0x16420,0x%h_0x%h\n0x16440,0x%h_0x%h\n0x16460,0x%h_0x%h\n0x16480,0x%h_0x%h\n0x164A0,0x%h_0x%h\n0x164C0,0x%h_0x%h\n0x164E0,0x%h_0x%h\n0x16500,0x%h_0x%h\n0x16520,0x%h_0x%h\n0x16540,0x%h_0x%h\n0x16560,0x%h_0x%h\n0x16580,0x%h_0x%h\n0x165A0,0x%h_0x%h\n0x165C0,0x%h_0x%h\n0x165E0,0x%h_0x%h\n0x16600,0x%h_0x%h\n0x16620,0x%h_0x%h\n0x16640,0x%h_0x%h\n0x16660,0x%h_0x%h\n0x16680,0x%h_0x%h\n0x166A0,0x%h_0x%h\n0x166C0,0x%h_0x%h\n0x166E0,0x%h_0x%h\n0x16700,0x%h_0x%h\n0x16720,0x%h_0x%h\n0x16740,0x%h_0x%h\n0x16760,0x%h_0x%h\n0x16780,0x%h_0x%h\n0x167A0,0x%h_0x%h\n0x167C0,0x%h_0x%h\n0x167E0,0x%h_0x%h\n0x16800,0x%h_0x%h\n0x16820,0x%h_0x%h\n0x16840,0x%h_0x%h\n0x16860,0x%h_0x%h\n0x16880,0x%h_0x%h\n0x168A0,0x%h_0x%h\n0x168C0,0x%h_0x%h\n0x168E0,0x%h_0x%h\n0x16900,0x%h_0x%h\n0x16920,0x%h_0x%h\n0x16940,0x%h_0x%h\n0x16960,0x%h_0x%h\n0x16980,0x%h_0x%h\n0x169A0,0x%h_0x%h\n0x169C0,0x%h_0x%h\n0x169E0,0x%h_0x%h\n0x16A00,0x%h_0x%h\n0x16A20,0x%h_0x%h\n0x16A40,0x%h_0x%h\n0x16A60,0x%h_0x%h\n0x16A80,0x%h_0x%h\n0x16AA0,0x%h_0x%h\n0x16AC0,0x%h_0x%h\n0x16AE0,0x%h_0x%h\n0x16B00,0x%h_0x%h\n0x16B20,0x%h_0x%h\n0x16B40,0x%h_0x%h\n0x16B60,0x%h_0x%h\n0x16B80,0x%h_0x%h\n0x16BA0,0x%h_0x%h\n0x16BC0,0x%h_0x%h\n0x16BE0,0x%h_0x%h\n0x16C00,0x%h_0x%h\n0x16C20,0x%h_0x%h\n0x16C40,0x%h_0x%h\n0x16C60,0x%h_0x%h\n0x16C80,0x%h_0x%h\n0x16CA0,0x%h_0x%h\n0x16CC0,0x%h_0x%h\n0x16CE0,0x%h_0x%h\n0x16D00,0x%h_0x%h\n0x16D20,0x%h_0x%h\n0x16D40,0x%h_0x%h\n0x16D60,0x%h_0x%h\n0x16D80,0x%h_0x%h\n0x16DA0,0x%h_0x%h\n0x16DC0,0x%h_0x%h\n0x16DE0,0x%h_0x%h\n0x16E00,0x%h_0x%h\n0x16E20,0x%h_0x%h\n0x16E40,0x%h_0x%h\n0x16E60,0x%h_0x%h\n0x16E80,0x%h_0x%h\n0x16EA0,0x%h_0x%h\n0x16EC0,0x%h_0x%h\n0x16EE0,0x%h_0x%h\n0x16F00,0x%h_0x%h\n0x16F20,0x%h_0x%h\n0x16F40,0x%h_0x%h\n0x16F60,0x%h_0x%h\n0x16F80,0x%h_0x%h\n0x16FA0,0x%h_0x%h\n0x16FC0,0x%h_0x%h\n0x16FE0,0x%h_0x%h\n0x17000,0x%h_0x%h\n0x17020,0x%h_0x%h\n0x17040,0x%h_0x%h\n0x17060,0x%h_0x%h\n0x17080,0x%h_0x%h\n0x170A0,0x%h_0x%h\n0x170C0,0x%h_0x%h\n0x170E0,0x%h_0x%h\n0x17100,0x%h_0x%h\n0x17120,0x%h_0x%h\n0x17140,0x%h_0x%h\n0x17160,0x%h_0x%h\n0x17180,0x%h_0x%h\n0x171A0,0x%h_0x%h\n0x171C0,0x%h_0x%h\n0x171E0,0x%h_0x%h\n0x17200,0x%h_0x%h\n0x17220,0x%h_0x%h\n0x17240,0x%h_0x%h\n0x17260,0x%h_0x%h\n0x17280,0x%h_0x%h\n0x172A0,0x%h_0x%h\n0x172C0,0x%h_0x%h\n0x172E0,0x%h_0x%h\n0x17300,0x%h_0x%h\n0x17320,0x%h_0x%h\n0x17340,0x%h_0x%h\n0x17360,0x%h_0x%h\n0x17380,0x%h_0x%h\n0x173A0,0x%h_0x%h\n0x173C0,0x%h_0x%h\n0x173E0,0x%h_0x%h\n0x17400,0x%h_0x%h\n0x17420,0x%h_0x%h\n0x17440,0x%h_0x%h\n0x17460,0x%h_0x%h\n0x17480,0x%h_0x%h\n0x174A0,0x%h_0x%h\n0x174C0,0x%h_0x%h\n0x174E0,0x%h_0x%h\n0x17500,0x%h_0x%h\n0x17520,0x%h_0x%h\n0x17540,0x%h_0x%h\n0x17560,0x%h_0x%h\n0x17580,0x%h_0x%h\n0x175A0,0x%h_0x%h\n0x175C0,0x%h_0x%h\n0x175E0,0x%h_0x%h\n0x17600,0x%h_0x%h\n0x17620,0x%h_0x%h\n0x17640,0x%h_0x%h\n0x17660,0x%h_0x%h\n0x17680,0x%h_0x%h\n0x176A0,0x%h_0x%h\n0x176C0,0x%h_0x%h\n0x176E0,0x%h_0x%h\n0x17700,0x%h_0x%h\n0x17720,0x%h_0x%h\n0x17740,0x%h_0x%h\n0x17760,0x%h_0x%h\n0x17780,0x%h_0x%h\n0x177A0,0x%h_0x%h\n0x177C0,0x%h_0x%h\n0x177E0,0x%h_0x%h\n0x17800,0x%h_0x%h\n0x17820,0x%h_0x%h\n0x17840,0x%h_0x%h\n0x17860,0x%h_0x%h\n0x17880,0x%h_0x%h\n0x178A0,0x%h_0x%h\n0x178C0,0x%h_0x%h\n0x178E0,0x%h_0x%h\n0x17900,0x%h_0x%h\n0x17920,0x%h_0x%h\n0x17940,0x%h_0x%h\n0x17960,0x%h_0x%h\n0x17980,0x%h_0x%h\n0x179A0,0x%h_0x%h\n0x179C0,0x%h_0x%h\n0x179E0,0x%h_0x%h\n0x17A00,0x%h_0x%h\n0x17A20,0x%h_0x%h\n0x17A40,0x%h_0x%h\n0x17A60,0x%h_0x%h\n0x17A80,0x%h_0x%h\n0x17AA0,0x%h_0x%h\n0x17AC0,0x%h_0x%h\n0x17AE0,0x%h_0x%h\n0x17B00,0x%h_0x%h\n0x17B20,0x%h_0x%h\n0x17B40,0x%h_0x%h\n0x17B60,0x%h_0x%h\n0x17B80,0x%h_0x%h\n0x17BA0,0x%h_0x%h\n0x17BC0,0x%h_0x%h\n0x17BE0,0x%h_0x%h\n0x17C00,0x%h_0x%h\n0x17C20,0x%h_0x%h\n0x17C40,0x%h_0x%h\n0x17C60,0x%h_0x%h\n0x17C80,0x%h_0x%h\n0x17CA0,0x%h_0x%h\n0x17CC0,0x%h_0x%h\n0x17CE0,0x%h_0x%h\n0x17D00,0x%h_0x%h\n0x17D20,0x%h_0x%h\n0x17D40,0x%h_0x%h\n0x17D60,0x%h_0x%h\n0x17D80,0x%h_0x%h\n0x17DA0,0x%h_0x%h\n0x17DC0,0x%h_0x%h\n0x17DE0,0x%h_0x%h\n0x17E00,0x%h_0x%h\n0x17E20,0x%h_0x%h\n0x17E40,0x%h_0x%h\n0x17E60,0x%h_0x%h\n0x17E80,0x%h_0x%h\n0x17EA0,0x%h_0x%h\n0x17EC0,0x%h_0x%h\n0x17EE0,0x%h_0x%h\n0x17F00,0x%h_0x%h\n0x17F20,0x%h_0x%h\n0x17F40,0x%h_0x%h\n0x17F60,0x%h_0x%h\n0x17F80,0x%h_0x%h\n0x17FA0,0x%h_0x%h\n0x17FC0,0x%h_0x%h\n0x17FE0,0x%h_0x%h\n0x18000,0x%h_0x%h\n0x18020,0x%h_0x%h\n0x18040,0x%h_0x%h\n0x18060,0x%h_0x%h\n0x18080,0x%h_0x%h\n0x180A0,0x%h_0x%h\n0x180C0,0x%h_0x%h\n0x180E0,0x%h_0x%h\n0x18100,0x%h_0x%h\n0x18120,0x%h_0x%h\n0x18140,0x%h_0x%h\n0x18160,0x%h_0x%h\n0x18180,0x%h_0x%h\n0x181A0,0x%h_0x%h\n0x181C0,0x%h_0x%h\n0x181E0,0x%h_0x%h\n0x18200,0x%h_0x%h\n0x18220,0x%h_0x%h\n0x18240,0x%h_0x%h\n0x18260,0x%h_0x%h\n0x18280,0x%h_0x%h\n0x182A0,0x%h_0x%h\n0x182C0,0x%h_0x%h\n0x182E0,0x%h_0x%h\n0x18300,0x%h_0x%h\n0x18320,0x%h_0x%h\n0x18340,0x%h_0x%h\n0x18360,0x%h_0x%h\n0x18380,0x%h_0x%h\n0x183A0,0x%h_0x%h\n0x183C0,0x%h_0x%h\n0x183E0,0x%h_0x%h\n0x18400,0x%h_0x%h\n0x18420,0x%h_0x%h\n0x18440,0x%h_0x%h\n0x18460,0x%h_0x%h\n0x18480,0x%h_0x%h\n0x184A0,0x%h_0x%h\n0x184C0,0x%h_0x%h\n0x184E0,0x%h_0x%h\n0x18500,0x%h_0x%h\n0x18520,0x%h_0x%h\n0x18540,0x%h_0x%h\n0x18560,0x%h_0x%h\n0x18580,0x%h_0x%h\n0x185A0,0x%h_0x%h\n0x185C0,0x%h_0x%h\n0x185E0,0x%h_0x%h\n0x18600,0x%h_0x%h\n0x18620,0x%h_0x%h\n0x18640,0x%h_0x%h\n0x18660,0x%h_0x%h\n0x18680,0x%h_0x%h\n0x186A0,0x%h_0x%h\n0x186C0,0x%h_0x%h\n0x186E0,0x%h_0x%h\n0x18700,0x%h_0x%h\n0x18720,0x%h_0x%h\n0x18740,0x%h_0x%h\n0x18760,0x%h_0x%h\n0x18780,0x%h_0x%h\n0x187A0,0x%h_0x%h\n0x187C0,0x%h_0x%h\n0x187E0,0x%h_0x%h\n0x18800,0x%h_0x%h\n0x18820,0x%h_0x%h\n0x18840,0x%h_0x%h\n0x18860,0x%h_0x%h\n0x18880,0x%h_0x%h\n0x188A0,0x%h_0x%h\n0x188C0,0x%h_0x%h\n0x188E0,0x%h_0x%h\n0x18900,0x%h_0x%h\n0x18920,0x%h_0x%h\n0x18940,0x%h_0x%h\n0x18960,0x%h_0x%h\n0x18980,0x%h_0x%h\n0x189A0,0x%h_0x%h\n0x189C0,0x%h_0x%h\n0x189E0,0x%h_0x%h\n0x18A00,0x%h_0x%h\n0x18A20,0x%h_0x%h\n0x18A40,0x%h_0x%h\n0x18A60,0x%h_0x%h\n0x18A80,0x%h_0x%h\n0x18AA0,0x%h_0x%h\n0x18AC0,0x%h_0x%h\n0x18AE0,0x%h_0x%h\n0x18B00,0x%h_0x%h\n0x18B20,0x%h_0x%h\n0x18B40,0x%h_0x%h\n0x18B60,0x%h_0x%h\n0x18B80,0x%h_0x%h\n0x18BA0,0x%h_0x%h\n0x18BC0,0x%h_0x%h\n0x18BE0,0x%h_0x%h\n0x18C00,0x%h_0x%h\n0x18C20,0x%h_0x%h\n0x18C40,0x%h_0x%h\n0x18C60,0x%h_0x%h\n0x18C80,0x%h_0x%h\n0x18CA0,0x%h_0x%h\n0x18CC0,0x%h_0x%h\n0x18CE0,0x%h_0x%h\n0x18D00,0x%h_0x%h\n0x18D20,0x%h_0x%h\n0x18D40,0x%h_0x%h\n0x18D60,0x%h_0x%h\n0x18D80,0x%h_0x%h\n0x18DA0,0x%h_0x%h\n0x18DC0,0x%h_0x%h\n0x18DE0,0x%h_0x%h\n0x18E00,0x%h_0x%h\n0x18E20,0x%h_0x%h\n0x18E40,0x%h_0x%h\n0x18E60,0x%h_0x%h\n0x18E80,0x%h_0x%h\n0x18EA0,0x%h_0x%h\n0x18EC0,0x%h_0x%h\n0x18EE0,0x%h_0x%h\n0x18F00,0x%h_0x%h\n0x18F20,0x%h_0x%h\n0x18F40,0x%h_0x%h\n0x18F60,0x%h_0x%h\n0x18F80,0x%h_0x%h\n0x18FA0,0x%h_0x%h\n0x18FC0,0x%h_0x%h\n0x18FE0,0x%h_0x%h\n0x19000,0x%h_0x%h\n0x19020,0x%h_0x%h\n0x19040,0x%h_0x%h\n0x19060,0x%h_0x%h\n0x19080,0x%h_0x%h\n0x190A0,0x%h_0x%h\n0x190C0,0x%h_0x%h\n0x190E0,0x%h_0x%h\n0x19100,0x%h_0x%h\n0x19120,0x%h_0x%h\n0x19140,0x%h_0x%h\n0x19160,0x%h_0x%h\n0x19180,0x%h_0x%h\n0x191A0,0x%h_0x%h\n0x191C0,0x%h_0x%h\n0x191E0,0x%h_0x%h\n0x19200,0x%h_0x%h\n0x19220,0x%h_0x%h\n0x19240,0x%h_0x%h\n0x19260,0x%h_0x%h\n0x19280,0x%h_0x%h\n0x192A0,0x%h_0x%h\n0x192C0,0x%h_0x%h\n0x192E0,0x%h_0x%h\n0x19300,0x%h_0x%h\n0x19320,0x%h_0x%h\n0x19340,0x%h_0x%h\n0x19360,0x%h_0x%h\n0x19380,0x%h_0x%h\n0x193A0,0x%h_0x%h\n0x193C0,0x%h_0x%h\n0x193E0,0x%h_0x%h\n0x19400,0x%h_0x%h\n0x19420,0x%h_0x%h\n0x19440,0x%h_0x%h\n0x19460,0x%h_0x%h\n0x19480,0x%h_0x%h\n0x194A0,0x%h_0x%h\n0x194C0,0x%h_0x%h\n0x194E0,0x%h_0x%h\n0x19500,0x%h_0x%h\n0x19520,0x%h_0x%h\n0x19540,0x%h_0x%h\n0x19560,0x%h_0x%h\n0x19580,0x%h_0x%h\n0x195A0,0x%h_0x%h\n0x195C0,0x%h_0x%h\n0x195E0,0x%h_0x%h\n0x19600,0x%h_0x%h\n0x19620,0x%h_0x%h\n0x19640,0x%h_0x%h\n0x19660,0x%h_0x%h\n0x19680,0x%h_0x%h\n0x196A0,0x%h_0x%h\n0x196C0,0x%h_0x%h\n0x196E0,0x%h_0x%h\n0x19700,0x%h_0x%h\n0x19720,0x%h_0x%h\n0x19740,0x%h_0x%h\n0x19760,0x%h_0x%h\n0x19780,0x%h_0x%h\n0x197A0,0x%h_0x%h\n0x197C0,0x%h_0x%h\n0x197E0,0x%h_0x%h\n0x19800,0x%h_0x%h\n0x19820,0x%h_0x%h\n0x19840,0x%h_0x%h\n0x19860,0x%h_0x%h\n0x19880,0x%h_0x%h\n0x198A0,0x%h_0x%h\n0x198C0,0x%h_0x%h\n0x198E0,0x%h_0x%h\n0x19900,0x%h_0x%h\n0x19920,0x%h_0x%h\n0x19940,0x%h_0x%h\n0x19960,0x%h_0x%h\n0x19980,0x%h_0x%h\n0x199A0,0x%h_0x%h\n0x199C0,0x%h_0x%h\n0x199E0,0x%h_0x%h\n0x19A00,0x%h_0x%h\n0x19A20,0x%h_0x%h\n0x19A40,0x%h_0x%h\n0x19A60,0x%h_0x%h\n0x19A80,0x%h_0x%h\n0x19AA0,0x%h_0x%h\n0x19AC0,0x%h_0x%h\n0x19AE0,0x%h_0x%h\n0x19B00,0x%h_0x%h\n0x19B20,0x%h_0x%h\n0x19B40,0x%h_0x%h\n0x19B60,0x%h_0x%h\n0x19B80,0x%h_0x%h\n0x19BA0,0x%h_0x%h\n0x19BC0,0x%h_0x%h\n0x19BE0,0x%h_0x%h\n0x19C00,0x%h_0x%h\n0x19C20,0x%h_0x%h\n0x19C40,0x%h_0x%h\n0x19C60,0x%h_0x%h\n0x19C80,0x%h_0x%h\n0x19CA0,0x%h_0x%h\n0x19CC0,0x%h_0x%h\n0x19CE0,0x%h_0x%h\n0x19D00,0x%h_0x%h\n0x19D20,0x%h_0x%h\n0x19D40,0x%h_0x%h\n0x19D60,0x%h_0x%h\n0x19D80,0x%h_0x%h\n0x19DA0,0x%h_0x%h\n0x19DC0,0x%h_0x%h\n0x19DE0,0x%h_0x%h\n0x19E00,0x%h_0x%h\n0x19E20,0x%h_0x%h\n0x19E40,0x%h_0x%h\n0x19E60,0x%h_0x%h\n0x19E80,0x%h_0x%h\n0x19EA0,0x%h_0x%h\n0x19EC0,0x%h_0x%h\n0x19EE0,0x%h_0x%h\n0x19F00,0x%h_0x%h\n0x19F20,0x%h_0x%h\n0x19F40,0x%h_0x%h\n0x19F60,0x%h_0x%h\n0x19F80,0x%h_0x%h\n0x19FA0,0x%h_0x%h\n0x19FC0,0x%h_0x%h\n0x19FE0,0x%h_0x%h\n0x1A000,0x%h_0x%h\n0x1A020,0x%h_0x%h\n0x1A040,0x%h_0x%h\n0x1A060,0x%h_0x%h\n0x1A080,0x%h_0x%h\n0x1A0A0,0x%h_0x%h\n0x1A0C0,0x%h_0x%h\n0x1A0E0,0x%h_0x%h\n0x1A100,0x%h_0x%h\n0x1A120,0x%h_0x%h\n0x1A140,0x%h_0x%h\n0x1A160,0x%h_0x%h\n0x1A180,0x%h_0x%h\n0x1A1A0,0x%h_0x%h\n0x1A1C0,0x%h_0x%h\n0x1A1E0,0x%h_0x%h\n0x1A200,0x%h_0x%h\n0x1A220,0x%h_0x%h\n0x1A240,0x%h_0x%h\n0x1A260,0x%h_0x%h\n0x1A280,0x%h_0x%h\n0x1A2A0,0x%h_0x%h\n0x1A2C0,0x%h_0x%h\n0x1A2E0,0x%h_0x%h\n0x1A300,0x%h_0x%h\n0x1A320,0x%h_0x%h\n0x1A340,0x%h_0x%h\n0x1A360,0x%h_0x%h\n0x1A380,0x%h_0x%h\n0x1A3A0,0x%h_0x%h\n0x1A3C0,0x%h_0x%h\n0x1A3E0,0x%h_0x%h\n0x1A400,0x%h_0x%h\n0x1A420,0x%h_0x%h\n0x1A440,0x%h_0x%h\n0x1A460,0x%h_0x%h\n0x1A480,0x%h_0x%h\n0x1A4A0,0x%h_0x%h\n0x1A4C0,0x%h_0x%h\n0x1A4E0,0x%h_0x%h\n0x1A500,0x%h_0x%h\n0x1A520,0x%h_0x%h\n0x1A540,0x%h_0x%h\n0x1A560,0x%h_0x%h\n0x1A580,0x%h_0x%h\n0x1A5A0,0x%h_0x%h\n0x1A5C0,0x%h_0x%h\n0x1A5E0,0x%h_0x%h\n0x1A600,0x%h_0x%h\n0x1A620,0x%h_0x%h\n0x1A640,0x%h_0x%h\n0x1A660,0x%h_0x%h\n0x1A680,0x%h_0x%h\n0x1A6A0,0x%h_0x%h\n0x1A6C0,0x%h_0x%h\n0x1A6E0,0x%h_0x%h\n0x1A700,0x%h_0x%h\n0x1A720,0x%h_0x%h\n0x1A740,0x%h_0x%h\n0x1A760,0x%h_0x%h\n0x1A780,0x%h_0x%h\n0x1A7A0,0x%h_0x%h\n0x1A7C0,0x%h_0x%h\n0x1A7E0,0x%h_0x%h\n0x1A800,0x%h_0x%h\n0x1A820,0x%h_0x%h\n0x1A840,0x%h_0x%h\n0x1A860,0x%h_0x%h\n0x1A880,0x%h_0x%h\n0x1A8A0,0x%h_0x%h\n0x1A8C0,0x%h_0x%h\n0x1A8E0,0x%h_0x%h\n0x1A900,0x%h_0x%h\n0x1A920,0x%h_0x%h\n0x1A940,0x%h_0x%h\n0x1A960,0x%h_0x%h\n0x1A980,0x%h_0x%h\n0x1A9A0,0x%h_0x%h\n0x1A9C0,0x%h_0x%h\n0x1A9E0,0x%h_0x%h\n0x1AA00,0x%h_0x%h\n0x1AA20,0x%h_0x%h\n0x1AA40,0x%h_0x%h\n0x1AA60,0x%h_0x%h\n0x1AA80,0x%h_0x%h\n0x1AAA0,0x%h_0x%h\n0x1AAC0,0x%h_0x%h\n0x1AAE0,0x%h_0x%h\n0x1AB00,0x%h_0x%h\n0x1AB20,0x%h_0x%h\n0x1AB40,0x%h_0x%h\n0x1AB60,0x%h_0x%h\n0x1AB80,0x%h_0x%h\n0x1ABA0,0x%h_0x%h\n0x1ABC0,0x%h_0x%h\n0x1ABE0,0x%h_0x%h\n0x1AC00,0x%h_0x%h\n0x1AC20,0x%h_0x%h\n0x1AC40,0x%h_0x%h\n0x1AC60,0x%h_0x%h\n0x1AC80,0x%h_0x%h\n0x1ACA0,0x%h_0x%h\n0x1ACC0,0x%h_0x%h\n0x1ACE0,0x%h_0x%h\n0x1AD00,0x%h_0x%h\n0x1AD20,0x%h_0x%h\n0x1AD40,0x%h_0x%h\n0x1AD60,0x%h_0x%h\n0x1AD80,0x%h_0x%h\n0x1ADA0,0x%h_0x%h\n0x1ADC0,0x%h_0x%h\n0x1ADE0,0x%h_0x%h\n0x1AE00,0x%h_0x%h\n0x1AE20,0x%h_0x%h\n0x1AE40,0x%h_0x%h\n0x1AE60,0x%h_0x%h\n0x1AE80,0x%h_0x%h\n0x1AEA0,0x%h_0x%h\n0x1AEC0,0x%h_0x%h\n0x1AEE0,0x%h_0x%h\n0x1AF00,0x%h_0x%h\n0x1AF20,0x%h_0x%h\n0x1AF40,0x%h_0x%h\n0x1AF60,0x%h_0x%h\n0x1AF80,0x%h_0x%h\n0x1AFA0,0x%h_0x%h\n0x1AFC0,0x%h_0x%h\n0x1AFE0,0x%h_0x%h\n0x1B000,0x%h_0x%h\n0x1B020,0x%h_0x%h\n0x1B040,0x%h_0x%h\n0x1B060,0x%h_0x%h\n0x1B080,0x%h_0x%h\n0x1B0A0,0x%h_0x%h\n0x1B0C0,0x%h_0x%h\n0x1B0E0,0x%h_0x%h\n0x1B100,0x%h_0x%h\n0x1B120,0x%h_0x%h\n0x1B140,0x%h_0x%h\n0x1B160,0x%h_0x%h\n0x1B180,0x%h_0x%h\n0x1B1A0,0x%h_0x%h\n0x1B1C0,0x%h_0x%h\n0x1B1E0,0x%h_0x%h\n0x1B200,0x%h_0x%h\n0x1B220,0x%h_0x%h\n0x1B240,0x%h_0x%h\n0x1B260,0x%h_0x%h\n0x1B280,0x%h_0x%h\n0x1B2A0,0x%h_0x%h\n0x1B2C0,0x%h_0x%h\n0x1B2E0,0x%h_0x%h\n0x1B300,0x%h_0x%h\n0x1B320,0x%h_0x%h\n0x1B340,0x%h_0x%h\n0x1B360,0x%h_0x%h\n0x1B380,0x%h_0x%h\n0x1B3A0,0x%h_0x%h\n0x1B3C0,0x%h_0x%h\n0x1B3E0,0x%h_0x%h\n0x1B400,0x%h_0x%h\n0x1B420,0x%h_0x%h\n0x1B440,0x%h_0x%h\n0x1B460,0x%h_0x%h\n0x1B480,0x%h_0x%h\n0x1B4A0,0x%h_0x%h\n0x1B4C0,0x%h_0x%h\n0x1B4E0,0x%h_0x%h\n0x1B500,0x%h_0x%h\n0x1B520,0x%h_0x%h\n0x1B540,0x%h_0x%h\n0x1B560,0x%h_0x%h\n0x1B580,0x%h_0x%h\n0x1B5A0,0x%h_0x%h\n0x1B5C0,0x%h_0x%h\n0x1B5E0,0x%h_0x%h\n0x1B600,0x%h_0x%h\n0x1B620,0x%h_0x%h\n0x1B640,0x%h_0x%h\n0x1B660,0x%h_0x%h\n0x1B680,0x%h_0x%h\n0x1B6A0,0x%h_0x%h\n0x1B6C0,0x%h_0x%h\n0x1B6E0,0x%h_0x%h\n0x1B700,0x%h_0x%h\n0x1B720,0x%h_0x%h\n0x1B740,0x%h_0x%h\n0x1B760,0x%h_0x%h\n0x1B780,0x%h_0x%h\n0x1B7A0,0x%h_0x%h\n0x1B7C0,0x%h_0x%h\n0x1B7E0,0x%h_0x%h\n0x1B800,0x%h_0x%h\n0x1B820,0x%h_0x%h\n0x1B840,0x%h_0x%h\n0x1B860,0x%h_0x%h\n0x1B880,0x%h_0x%h\n0x1B8A0,0x%h_0x%h\n0x1B8C0,0x%h_0x%h\n0x1B8E0,0x%h_0x%h\n0x1B900,0x%h_0x%h\n0x1B920,0x%h_0x%h\n0x1B940,0x%h_0x%h\n0x1B960,0x%h_0x%h\n0x1B980,0x%h_0x%h\n0x1B9A0,0x%h_0x%h\n0x1B9C0,0x%h_0x%h\n0x1B9E0,0x%h_0x%h\n0x1BA00,0x%h_0x%h\n0x1BA20,0x%h_0x%h\n0x1BA40,0x%h_0x%h\n0x1BA60,0x%h_0x%h\n0x1BA80,0x%h_0x%h\n0x1BAA0,0x%h_0x%h\n0x1BAC0,0x%h_0x%h\n0x1BAE0,0x%h_0x%h\n0x1BB00,0x%h_0x%h\n0x1BB20,0x%h_0x%h\n0x1BB40,0x%h_0x%h\n0x1BB60,0x%h_0x%h\n0x1BB80,0x%h_0x%h\n0x1BBA0,0x%h_0x%h\n0x1BBC0,0x%h_0x%h\n0x1BBE0,0x%h_0x%h\n0x1BC00,0x%h_0x%h\n0x1BC20,0x%h_0x%h\n0x1BC40,0x%h_0x%h\n0x1BC60,0x%h_0x%h\n0x1BC80,0x%h_0x%h\n0x1BCA0,0x%h_0x%h\n0x1BCC0,0x%h_0x%h\n0x1BCE0,0x%h_0x%h\n0x1BD00,0x%h_0x%h\n0x1BD20,0x%h_0x%h\n0x1BD40,0x%h_0x%h\n0x1BD60,0x%h_0x%h\n0x1BD80,0x%h_0x%h\n0x1BDA0,0x%h_0x%h\n0x1BDC0,0x%h_0x%h\n0x1BDE0,0x%h_0x%h\n0x1BE00,0x%h_0x%h\n0x1BE20,0x%h_0x%h\n0x1BE40,0x%h_0x%h\n0x1BE60,0x%h_0x%h\n0x1BE80,0x%h_0x%h\n0x1BEA0,0x%h_0x%h\n0x1BEC0,0x%h_0x%h\n0x1BEE0,0x%h_0x%h\n0x1BF00,0x%h_0x%h\n0x1BF20,0x%h_0x%h\n0x1BF40,0x%h_0x%h\n0x1BF60,0x%h_0x%h\n0x1BF80,0x%h_0x%h\n0x1BFA0,0x%h_0x%h\n0x1BFC0,0x%h_0x%h\n0x1BFE0,0x%h_0x%h\n0x1C000,0x%h_0x%h\n0x1C020,0x%h_0x%h\n0x1C040,0x%h_0x%h\n0x1C060,0x%h_0x%h\n0x1C080,0x%h_0x%h\n0x1C0A0,0x%h_0x%h\n0x1C0C0,0x%h_0x%h\n0x1C0E0,0x%h_0x%h\n0x1C100,0x%h_0x%h\n0x1C120,0x%h_0x%h\n0x1C140,0x%h_0x%h\n0x1C160,0x%h_0x%h\n0x1C180,0x%h_0x%h\n0x1C1A0,0x%h_0x%h\n0x1C1C0,0x%h_0x%h\n0x1C1E0,0x%h_0x%h\n0x1C200,0x%h_0x%h\n0x1C220,0x%h_0x%h\n0x1C240,0x%h_0x%h\n0x1C260,0x%h_0x%h\n0x1C280,0x%h_0x%h\n0x1C2A0,0x%h_0x%h\n0x1C2C0,0x%h_0x%h\n0x1C2E0,0x%h_0x%h\n0x1C300,0x%h_0x%h\n0x1C320,0x%h_0x%h\n0x1C340,0x%h_0x%h\n0x1C360,0x%h_0x%h\n0x1C380,0x%h_0x%h\n0x1C3A0,0x%h_0x%h\n0x1C3C0,0x%h_0x%h\n0x1C3E0,0x%h_0x%h\n0x1C400,0x%h_0x%h\n0x1C420,0x%h_0x%h\n0x1C440,0x%h_0x%h\n0x1C460,0x%h_0x%h\n0x1C480,0x%h_0x%h\n0x1C4A0,0x%h_0x%h\n0x1C4C0,0x%h_0x%h\n0x1C4E0,0x%h_0x%h\n0x1C500,0x%h_0x%h\n0x1C520,0x%h_0x%h\n0x1C540,0x%h_0x%h\n0x1C560,0x%h_0x%h\n0x1C580,0x%h_0x%h\n0x1C5A0,0x%h_0x%h\n0x1C5C0,0x%h_0x%h\n0x1C5E0,0x%h_0x%h\n0x1C600,0x%h_0x%h\n0x1C620,0x%h_0x%h\n0x1C640,0x%h_0x%h\n0x1C660,0x%h_0x%h\n0x1C680,0x%h_0x%h\n0x1C6A0,0x%h_0x%h\n0x1C6C0,0x%h_0x%h\n0x1C6E0,0x%h_0x%h\n0x1C700,0x%h_0x%h\n0x1C720,0x%h_0x%h\n0x1C740,0x%h_0x%h\n0x1C760,0x%h_0x%h\n0x1C780,0x%h_0x%h\n0x1C7A0,0x%h_0x%h\n0x1C7C0,0x%h_0x%h\n0x1C7E0,0x%h_0x%h\n0x1C800,0x%h_0x%h\n0x1C820,0x%h_0x%h\n0x1C840,0x%h_0x%h\n0x1C860,0x%h_0x%h\n0x1C880,0x%h_0x%h\n0x1C8A0,0x%h_0x%h\n0x1C8C0,0x%h_0x%h\n0x1C8E0,0x%h_0x%h\n0x1C900,0x%h_0x%h\n0x1C920,0x%h_0x%h\n0x1C940,0x%h_0x%h\n0x1C960,0x%h_0x%h\n0x1C980,0x%h_0x%h\n0x1C9A0,0x%h_0x%h\n0x1C9C0,0x%h_0x%h\n0x1C9E0,0x%h_0x%h\n0x1CA00,0x%h_0x%h\n0x1CA20,0x%h_0x%h\n0x1CA40,0x%h_0x%h\n0x1CA60,0x%h_0x%h\n0x1CA80,0x%h_0x%h\n0x1CAA0,0x%h_0x%h\n0x1CAC0,0x%h_0x%h\n0x1CAE0,0x%h_0x%h\n0x1CB00,0x%h_0x%h\n0x1CB20,0x%h_0x%h\n0x1CB40,0x%h_0x%h\n0x1CB60,0x%h_0x%h\n0x1CB80,0x%h_0x%h\n0x1CBA0,0x%h_0x%h\n0x1CBC0,0x%h_0x%h\n0x1CBE0,0x%h_0x%h\n0x1CC00,0x%h_0x%h\n0x1CC20,0x%h_0x%h\n0x1CC40,0x%h_0x%h\n0x1CC60,0x%h_0x%h\n0x1CC80,0x%h_0x%h\n0x1CCA0,0x%h_0x%h\n0x1CCC0,0x%h_0x%h\n0x1CCE0,0x%h_0x%h\n0x1CD00,0x%h_0x%h\n0x1CD20,0x%h_0x%h\n0x1CD40,0x%h_0x%h\n0x1CD60,0x%h_0x%h\n0x1CD80,0x%h_0x%h\n0x1CDA0,0x%h_0x%h\n0x1CDC0,0x%h_0x%h\n0x1CDE0,0x%h_0x%h\n0x1CE00,0x%h_0x%h\n0x1CE20,0x%h_0x%h\n0x1CE40,0x%h_0x%h\n0x1CE60,0x%h_0x%h\n0x1CE80,0x%h_0x%h\n0x1CEA0,0x%h_0x%h\n0x1CEC0,0x%h_0x%h\n0x1CEE0,0x%h_0x%h\n0x1CF00,0x%h_0x%h\n0x1CF20,0x%h_0x%h\n0x1CF40,0x%h_0x%h\n0x1CF60,0x%h_0x%h\n0x1CF80,0x%h_0x%h\n0x1CFA0,0x%h_0x%h\n0x1CFC0,0x%h_0x%h\n0x1CFE0,0x%h_0x%h\n0x1D000,0x%h_0x%h\n0x1D020,0x%h_0x%h\n0x1D040,0x%h_0x%h\n0x1D060,0x%h_0x%h\n0x1D080,0x%h_0x%h\n0x1D0A0,0x%h_0x%h\n0x1D0C0,0x%h_0x%h\n0x1D0E0,0x%h_0x%h\n0x1D100,0x%h_0x%h\n0x1D120,0x%h_0x%h\n0x1D140,0x%h_0x%h\n0x1D160,0x%h_0x%h\n0x1D180,0x%h_0x%h\n0x1D1A0,0x%h_0x%h\n0x1D1C0,0x%h_0x%h\n0x1D1E0,0x%h_0x%h\n0x1D200,0x%h_0x%h\n0x1D220,0x%h_0x%h\n0x1D240,0x%h_0x%h\n0x1D260,0x%h_0x%h\n0x1D280,0x%h_0x%h\n0x1D2A0,0x%h_0x%h\n0x1D2C0,0x%h_0x%h\n0x1D2E0,0x%h_0x%h\n0x1D300,0x%h_0x%h\n0x1D320,0x%h_0x%h\n0x1D340,0x%h_0x%h\n0x1D360,0x%h_0x%h\n0x1D380,0x%h_0x%h\n0x1D3A0,0x%h_0x%h\n0x1D3C0,0x%h_0x%h\n0x1D3E0,0x%h_0x%h\n0x1D400,0x%h_0x%h\n0x1D420,0x%h_0x%h\n0x1D440,0x%h_0x%h\n0x1D460,0x%h_0x%h\n0x1D480,0x%h_0x%h\n0x1D4A0,0x%h_0x%h\n0x1D4C0,0x%h_0x%h\n0x1D4E0,0x%h_0x%h\n0x1D500,0x%h_0x%h\n0x1D520,0x%h_0x%h\n0x1D540,0x%h_0x%h\n0x1D560,0x%h_0x%h\n0x1D580,0x%h_0x%h\n0x1D5A0,0x%h_0x%h\n0x1D5C0,0x%h_0x%h\n0x1D5E0,0x%h_0x%h\n0x1D600,0x%h_0x%h\n0x1D620,0x%h_0x%h\n0x1D640,0x%h_0x%h\n0x1D660,0x%h_0x%h\n0x1D680,0x%h_0x%h\n0x1D6A0,0x%h_0x%h\n0x1D6C0,0x%h_0x%h\n0x1D6E0,0x%h_0x%h\n0x1D700,0x%h_0x%h\n0x1D720,0x%h_0x%h\n0x1D740,0x%h_0x%h\n0x1D760,0x%h_0x%h\n0x1D780,0x%h_0x%h\n0x1D7A0,0x%h_0x%h\n0x1D7C0,0x%h_0x%h\n0x1D7E0,0x%h_0x%h\n0x1D800,0x%h_0x%h\n0x1D820,0x%h_0x%h\n0x1D840,0x%h_0x%h\n0x1D860,0x%h_0x%h\n0x1D880,0x%h_0x%h\n0x1D8A0,0x%h_0x%h\n0x1D8C0,0x%h_0x%h\n0x1D8E0,0x%h_0x%h\n0x1D900,0x%h_0x%h\n0x1D920,0x%h_0x%h\n0x1D940,0x%h_0x%h\n0x1D960,0x%h_0x%h\n0x1D980,0x%h_0x%h\n0x1D9A0,0x%h_0x%h\n0x1D9C0,0x%h_0x%h\n0x1D9E0,0x%h_0x%h\n0x1DA00,0x%h_0x%h\n0x1DA20,0x%h_0x%h\n0x1DA40,0x%h_0x%h\n0x1DA60,0x%h_0x%h\n0x1DA80,0x%h_0x%h\n0x1DAA0,0x%h_0x%h\n0x1DAC0,0x%h_0x%h\n0x1DAE0,0x%h_0x%h\n0x1DB00,0x%h_0x%h\n0x1DB20,0x%h_0x%h\n0x1DB40,0x%h_0x%h\n0x1DB60,0x%h_0x%h\n0x1DB80,0x%h_0x%h\n0x1DBA0,0x%h_0x%h\n0x1DBC0,0x%h_0x%h\n0x1DBE0,0x%h_0x%h\n0x1DC00,0x%h_0x%h\n0x1DC20,0x%h_0x%h\n0x1DC40,0x%h_0x%h\n0x1DC60,0x%h_0x%h\n0x1DC80,0x%h_0x%h\n0x1DCA0,0x%h_0x%h\n0x1DCC0,0x%h_0x%h\n0x1DCE0,0x%h_0x%h\n0x1DD00,0x%h_0x%h\n0x1DD20,0x%h_0x%h\n0x1DD40,0x%h_0x%h\n0x1DD60,0x%h_0x%h\n0x1DD80,0x%h_0x%h\n0x1DDA0,0x%h_0x%h\n0x1DDC0,0x%h_0x%h\n0x1DDE0,0x%h_0x%h\n0x1DE00,0x%h_0x%h\n0x1DE20,0x%h_0x%h\n0x1DE40,0x%h_0x%h\n0x1DE60,0x%h_0x%h\n0x1DE80,0x%h_0x%h\n0x1DEA0,0x%h_0x%h\n0x1DEC0,0x%h_0x%h\n0x1DEE0,0x%h_0x%h\n0x1DF00,0x%h_0x%h\n0x1DF20,0x%h_0x%h\n0x1DF40,0x%h_0x%h\n0x1DF60,0x%h_0x%h\n0x1DF80,0x%h_0x%h\n0x1DFA0,0x%h_0x%h\n0x1DFC0,0x%h_0x%h\n0x1DFE0,0x%h_0x%h\n0x1E000,0x%h_0x%h\n0x1E020,0x%h_0x%h\n0x1E040,0x%h_0x%h\n0x1E060,0x%h_0x%h\n0x1E080,0x%h_0x%h\n0x1E0A0,0x%h_0x%h\n0x1E0C0,0x%h_0x%h\n0x1E0E0,0x%h_0x%h\n0x1E100,0x%h_0x%h\n0x1E120,0x%h_0x%h\n0x1E140,0x%h_0x%h\n0x1E160,0x%h_0x%h\n0x1E180,0x%h_0x%h\n0x1E1A0,0x%h_0x%h\n0x1E1C0,0x%h_0x%h\n0x1E1E0,0x%h_0x%h\n0x1E200,0x%h_0x%h\n0x1E220,0x%h_0x%h\n0x1E240,0x%h_0x%h\n0x1E260,0x%h_0x%h\n0x1E280,0x%h_0x%h\n0x1E2A0,0x%h_0x%h\n0x1E2C0,0x%h_0x%h\n0x1E2E0,0x%h_0x%h\n0x1E300,0x%h_0x%h\n0x1E320,0x%h_0x%h\n0x1E340,0x%h_0x%h\n0x1E360,0x%h_0x%h\n0x1E380,0x%h_0x%h\n0x1E3A0,0x%h_0x%h\n0x1E3C0,0x%h_0x%h\n0x1E3E0,0x%h_0x%h\n0x1E400,0x%h_0x%h\n0x1E420,0x%h_0x%h\n0x1E440,0x%h_0x%h\n0x1E460,0x%h_0x%h\n0x1E480,0x%h_0x%h\n0x1E4A0,0x%h_0x%h\n0x1E4C0,0x%h_0x%h\n0x1E4E0,0x%h_0x%h\n0x1E500,0x%h_0x%h\n0x1E520,0x%h_0x%h\n0x1E540,0x%h_0x%h\n0x1E560,0x%h_0x%h\n0x1E580,0x%h_0x%h\n0x1E5A0,0x%h_0x%h\n0x1E5C0,0x%h_0x%h\n0x1E5E0,0x%h_0x%h\n0x1E600,0x%h_0x%h\n0x1E620,0x%h_0x%h\n0x1E640,0x%h_0x%h\n0x1E660,0x%h_0x%h\n0x1E680,0x%h_0x%h\n0x1E6A0,0x%h_0x%h\n0x1E6C0,0x%h_0x%h\n0x1E6E0,0x%h_0x%h\n0x1E700,0x%h_0x%h\n0x1E720,0x%h_0x%h\n0x1E740,0x%h_0x%h\n0x1E760,0x%h_0x%h\n0x1E780,0x%h_0x%h\n0x1E7A0,0x%h_0x%h\n0x1E7C0,0x%h_0x%h\n0x1E7E0,0x%h_0x%h\n0x1E800,0x%h_0x%h\n0x1E820,0x%h_0x%h\n0x1E840,0x%h_0x%h\n0x1E860,0x%h_0x%h\n0x1E880,0x%h_0x%h\n0x1E8A0,0x%h_0x%h\n0x1E8C0,0x%h_0x%h\n0x1E8E0,0x%h_0x%h\n0x1E900,0x%h_0x%h\n0x1E920,0x%h_0x%h\n0x1E940,0x%h_0x%h\n0x1E960,0x%h_0x%h\n0x1E980,0x%h_0x%h\n0x1E9A0,0x%h_0x%h\n0x1E9C0,0x%h_0x%h\n0x1E9E0,0x%h_0x%h\n0x1EA00,0x%h_0x%h\n0x1EA20,0x%h_0x%h\n0x1EA40,0x%h_0x%h\n0x1EA60,0x%h_0x%h\n0x1EA80,0x%h_0x%h\n0x1EAA0,0x%h_0x%h\n0x1EAC0,0x%h_0x%h\n0x1EAE0,0x%h_0x%h\n0x1EB00,0x%h_0x%h\n0x1EB20,0x%h_0x%h\n0x1EB40,0x%h_0x%h\n0x1EB60,0x%h_0x%h\n0x1EB80,0x%h_0x%h\n0x1EBA0,0x%h_0x%h\n0x1EBC0,0x%h_0x%h\n0x1EBE0,0x%h_0x%h\n0x1EC00,0x%h_0x%h\n0x1EC20,0x%h_0x%h\n0x1EC40,0x%h_0x%h\n0x1EC60,0x%h_0x%h\n0x1EC80,0x%h_0x%h\n0x1ECA0,0x%h_0x%h\n0x1ECC0,0x%h_0x%h\n0x1ECE0,0x%h_0x%h\n0x1ED00,0x%h_0x%h\n0x1ED20,0x%h_0x%h\n0x1ED40,0x%h_0x%h\n0x1ED60,0x%h_0x%h\n0x1ED80,0x%h_0x%h\n0x1EDA0,0x%h_0x%h\n0x1EDC0,0x%h_0x%h\n0x1EDE0,0x%h_0x%h\n0x1EE00,0x%h_0x%h\n0x1EE20,0x%h_0x%h\n0x1EE40,0x%h_0x%h\n0x1EE60,0x%h_0x%h\n0x1EE80,0x%h_0x%h\n0x1EEA0,0x%h_0x%h\n0x1EEC0,0x%h_0x%h\n0x1EEE0,0x%h_0x%h\n0x1EF00,0x%h_0x%h\n0x1EF20,0x%h_0x%h\n0x1EF40,0x%h_0x%h\n0x1EF60,0x%h_0x%h\n0x1EF80,0x%h_0x%h\n0x1EFA0,0x%h_0x%h\n0x1EFC0,0x%h_0x%h\n0x1EFE0,0x%h_0x%h\n0x1F000,0x%h_0x%h\n0x1F020,0x%h_0x%h\n0x1F040,0x%h_0x%h\n0x1F060,0x%h_0x%h\n0x1F080,0x%h_0x%h\n0x1F0A0,0x%h_0x%h\n0x1F0C0,0x%h_0x%h\n0x1F0E0,0x%h_0x%h\n0x1F100,0x%h_0x%h\n0x1F120,0x%h_0x%h\n0x1F140,0x%h_0x%h\n0x1F160,0x%h_0x%h\n0x1F180,0x%h_0x%h\n0x1F1A0,0x%h_0x%h\n0x1F1C0,0x%h_0x%h\n0x1F1E0,0x%h_0x%h\n0x1F200,0x%h_0x%h\n0x1F220,0x%h_0x%h\n0x1F240,0x%h_0x%h\n0x1F260,0x%h_0x%h\n0x1F280,0x%h_0x%h\n0x1F2A0,0x%h_0x%h\n0x1F2C0,0x%h_0x%h\n0x1F2E0,0x%h_0x%h\n0x1F300,0x%h_0x%h\n0x1F320,0x%h_0x%h\n0x1F340,0x%h_0x%h\n0x1F360,0x%h_0x%h\n0x1F380,0x%h_0x%h\n0x1F3A0,0x%h_0x%h\n0x1F3C0,0x%h_0x%h\n0x1F3E0,0x%h_0x%h\n0x1F400,0x%h_0x%h\n0x1F420,0x%h_0x%h\n0x1F440,0x%h_0x%h\n0x1F460,0x%h_0x%h\n0x1F480,0x%h_0x%h\n0x1F4A0,0x%h_0x%h\n0x1F4C0,0x%h_0x%h\n0x1F4E0,0x%h_0x%h\n0x1F500,0x%h_0x%h\n0x1F520,0x%h_0x%h\n0x1F540,0x%h_0x%h\n0x1F560,0x%h_0x%h\n0x1F580,0x%h_0x%h\n0x1F5A0,0x%h_0x%h\n0x1F5C0,0x%h_0x%h\n0x1F5E0,0x%h_0x%h\n0x1F600,0x%h_0x%h\n0x1F620,0x%h_0x%h\n0x1F640,0x%h_0x%h\n0x1F660,0x%h_0x%h\n0x1F680,0x%h_0x%h\n0x1F6A0,0x%h_0x%h\n0x1F6C0,0x%h_0x%h\n0x1F6E0,0x%h_0x%h\n0x1F700,0x%h_0x%h\n0x1F720,0x%h_0x%h\n0x1F740,0x%h_0x%h\n0x1F760,0x%h_0x%h\n0x1F780,0x%h_0x%h\n0x1F7A0,0x%h_0x%h\n0x1F7C0,0x%h_0x%h\n0x1F7E0,0x%h_0x%h\n0x1F800,0x%h_0x%h\n0x1F820,0x%h_0x%h\n0x1F840,0x%h_0x%h\n0x1F860,0x%h_0x%h\n0x1F880,0x%h_0x%h\n0x1F8A0,0x%h_0x%h\n0x1F8C0,0x%h_0x%h\n0x1F8E0,0x%h_0x%h\n0x1F900,0x%h_0x%h\n0x1F920,0x%h_0x%h\n0x1F940,0x%h_0x%h\n0x1F960,0x%h_0x%h\n0x1F980,0x%h_0x%h\n0x1F9A0,0x%h_0x%h\n0x1F9C0,0x%h_0x%h\n0x1F9E0,0x%h_0x%h\n0x1FA00,0x%h_0x%h\n0x1FA20,0x%h_0x%h\n0x1FA40,0x%h_0x%h\n0x1FA60,0x%h_0x%h\n0x1FA80,0x%h_0x%h\n0x1FAA0,0x%h_0x%h\n0x1FAC0,0x%h_0x%h\n0x1FAE0,0x%h_0x%h\n0x1FB00,0x%h_0x%h\n0x1FB20,0x%h_0x%h\n0x1FB40,0x%h_0x%h\n0x1FB60,0x%h_0x%h\n0x1FB80,0x%h_0x%h\n0x1FBA0,0x%h_0x%h\n0x1FBC0,0x%h_0x%h\n0x1FBE0,0x%h_0x%h\n0x1FC00,0x%h_0x%h\n0x1FC20,0x%h_0x%h\n0x1FC40,0x%h_0x%h\n0x1FC60,0x%h_0x%h\n0x1FC80,0x%h_0x%h\n0x1FCA0,0x%h_0x%h\n0x1FCC0,0x%h_0x%h\n0x1FCE0,0x%h_0x%h\n0x1FD00,0x%h_0x%h\n0x1FD20,0x%h_0x%h\n0x1FD40,0x%h_0x%h\n0x1FD60,0x%h_0x%h\n0x1FD80,0x%h_0x%h\n0x1FDA0,0x%h_0x%h\n0x1FDC0,0x%h_0x%h\n0x1FDE0,0x%h_0x%h\n0x1FE00,0x%h_0x%h\n0x1FE20,0x%h_0x%h\n0x1FE40,0x%h_0x%h\n0x1FE60,0x%h_0x%h\n0x1FE80,0x%h_0x%h\n0x1FEA0,0x%h_0x%h\n0x1FEC0,0x%h_0x%h\n0x1FEE0,0x%h_0x%h\n0x1FF00,0x%h_0x%h\n0x1FF20,0x%h_0x%h\n0x1FF40,0x%h_0x%h\n0x1FF60,0x%h_0x%h\n0x1FF80,0x%h_0x%h\n0x1FFA0,0x%h_0x%h\n0x1FFC0,0x%h_0x%h\n0x1FFE0,0x%h_0x%h\n",db_odd.mem_bank[0],db_even.mem_bank[0],db_odd.mem_bank[1],db_even.mem_bank[1],db_odd.mem_bank[2],db_even.mem_bank[2],db_odd.mem_bank[3],db_even.mem_bank[3],db_odd.mem_bank[4],db_even.mem_bank[4],db_odd.mem_bank[5],db_even.mem_bank[5],db_odd.mem_bank[6],db_even.mem_bank[6],db_odd.mem_bank[7],db_even.mem_bank[7],db_odd.mem_bank[8],db_even.mem_bank[8],db_odd.mem_bank[9],db_even.mem_bank[9],db_odd.mem_bank[10],db_even.mem_bank[10],db_odd.mem_bank[11],db_even.mem_bank[11],db_odd.mem_bank[12],db_even.mem_bank[12],db_odd.mem_bank[13],db_even.mem_bank[13],db_odd.mem_bank[14],db_even.mem_bank[14],db_odd.mem_bank[15],db_even.mem_bank[15],db_odd.mem_bank[16],db_even.mem_bank[16],db_odd.mem_bank[17],db_even.mem_bank[17],db_odd.mem_bank[18],db_even.mem_bank[18],db_odd.mem_bank[19],db_even.mem_bank[19],db_odd.mem_bank[20],db_even.mem_bank[20],db_odd.mem_bank[21],db_even.mem_bank[21],db_odd.mem_bank[22],db_even.mem_bank[22],db_odd.mem_bank[23],db_even.mem_bank[23],db_odd.mem_bank[24],db_even.mem_bank[24],db_odd.mem_bank[25],db_even.mem_bank[25],db_odd.mem_bank[26],db_even.mem_bank[26],db_odd.mem_bank[27],db_even.mem_bank[27],db_odd.mem_bank[28],db_even.mem_bank[28],db_odd.mem_bank[29],db_even.mem_bank[29],db_odd.mem_bank[30],db_even.mem_bank[30],db_odd.mem_bank[31],db_even.mem_bank[31],db_odd.mem_bank[32],db_even.mem_bank[32],db_odd.mem_bank[33],db_even.mem_bank[33],db_odd.mem_bank[34],db_even.mem_bank[34],db_odd.mem_bank[35],db_even.mem_bank[35],db_odd.mem_bank[36],db_even.mem_bank[36],db_odd.mem_bank[37],db_even.mem_bank[37],db_odd.mem_bank[38],db_even.mem_bank[38],db_odd.mem_bank[39],db_even.mem_bank[39],db_odd.mem_bank[40],db_even.mem_bank[40],db_odd.mem_bank[41],db_even.mem_bank[41],db_odd.mem_bank[42],db_even.mem_bank[42],db_odd.mem_bank[43],db_even.mem_bank[43],db_odd.mem_bank[44],db_even.mem_bank[44],db_odd.mem_bank[45],db_even.mem_bank[45],db_odd.mem_bank[46],db_even.mem_bank[46],db_odd.mem_bank[47],db_even.mem_bank[47],db_odd.mem_bank[48],db_even.mem_bank[48],db_odd.mem_bank[49],db_even.mem_bank[49],db_odd.mem_bank[50],db_even.mem_bank[50],db_odd.mem_bank[51],db_even.mem_bank[51],db_odd.mem_bank[52],db_even.mem_bank[52],db_odd.mem_bank[53],db_even.mem_bank[53],db_odd.mem_bank[54],db_even.mem_bank[54],db_odd.mem_bank[55],db_even.mem_bank[55],db_odd.mem_bank[56],db_even.mem_bank[56],db_odd.mem_bank[57],db_even.mem_bank[57],db_odd.mem_bank[58],db_even.mem_bank[58],db_odd.mem_bank[59],db_even.mem_bank[59],db_odd.mem_bank[60],db_even.mem_bank[60],db_odd.mem_bank[61],db_even.mem_bank[61],db_odd.mem_bank[62],db_even.mem_bank[62],db_odd.mem_bank[63],db_even.mem_bank[63],db_odd.mem_bank[64],db_even.mem_bank[64],db_odd.mem_bank[65],db_even.mem_bank[65],db_odd.mem_bank[66],db_even.mem_bank[66],db_odd.mem_bank[67],db_even.mem_bank[67],db_odd.mem_bank[68],db_even.mem_bank[68],db_odd.mem_bank[69],db_even.mem_bank[69],db_odd.mem_bank[70],db_even.mem_bank[70],db_odd.mem_bank[71],db_even.mem_bank[71],db_odd.mem_bank[72],db_even.mem_bank[72],db_odd.mem_bank[73],db_even.mem_bank[73],db_odd.mem_bank[74],db_even.mem_bank[74],db_odd.mem_bank[75],db_even.mem_bank[75],db_odd.mem_bank[76],db_even.mem_bank[76],db_odd.mem_bank[77],db_even.mem_bank[77],db_odd.mem_bank[78],db_even.mem_bank[78],db_odd.mem_bank[79],db_even.mem_bank[79],db_odd.mem_bank[80],db_even.mem_bank[80],db_odd.mem_bank[81],db_even.mem_bank[81],db_odd.mem_bank[82],db_even.mem_bank[82],db_odd.mem_bank[83],db_even.mem_bank[83],db_odd.mem_bank[84],db_even.mem_bank[84],db_odd.mem_bank[85],db_even.mem_bank[85],db_odd.mem_bank[86],db_even.mem_bank[86],db_odd.mem_bank[87],db_even.mem_bank[87],db_odd.mem_bank[88],db_even.mem_bank[88],db_odd.mem_bank[89],db_even.mem_bank[89],db_odd.mem_bank[90],db_even.mem_bank[90],db_odd.mem_bank[91],db_even.mem_bank[91],db_odd.mem_bank[92],db_even.mem_bank[92],db_odd.mem_bank[93],db_even.mem_bank[93],db_odd.mem_bank[94],db_even.mem_bank[94],db_odd.mem_bank[95],db_even.mem_bank[95],db_odd.mem_bank[96],db_even.mem_bank[96],db_odd.mem_bank[97],db_even.mem_bank[97],db_odd.mem_bank[98],db_even.mem_bank[98],db_odd.mem_bank[99],db_even.mem_bank[99],db_odd.mem_bank[100],db_even.mem_bank[100],db_odd.mem_bank[101],db_even.mem_bank[101],db_odd.mem_bank[102],db_even.mem_bank[102],db_odd.mem_bank[103],db_even.mem_bank[103],db_odd.mem_bank[104],db_even.mem_bank[104],db_odd.mem_bank[105],db_even.mem_bank[105],db_odd.mem_bank[106],db_even.mem_bank[106],db_odd.mem_bank[107],db_even.mem_bank[107],db_odd.mem_bank[108],db_even.mem_bank[108],db_odd.mem_bank[109],db_even.mem_bank[109],db_odd.mem_bank[110],db_even.mem_bank[110],db_odd.mem_bank[111],db_even.mem_bank[111],db_odd.mem_bank[112],db_even.mem_bank[112],db_odd.mem_bank[113],db_even.mem_bank[113],db_odd.mem_bank[114],db_even.mem_bank[114],db_odd.mem_bank[115],db_even.mem_bank[115],db_odd.mem_bank[116],db_even.mem_bank[116],db_odd.mem_bank[117],db_even.mem_bank[117],db_odd.mem_bank[118],db_even.mem_bank[118],db_odd.mem_bank[119],db_even.mem_bank[119],db_odd.mem_bank[120],db_even.mem_bank[120],db_odd.mem_bank[121],db_even.mem_bank[121],db_odd.mem_bank[122],db_even.mem_bank[122],db_odd.mem_bank[123],db_even.mem_bank[123],db_odd.mem_bank[124],db_even.mem_bank[124],db_odd.mem_bank[125],db_even.mem_bank[125],db_odd.mem_bank[126],db_even.mem_bank[126],db_odd.mem_bank[127],db_even.mem_bank[127],db_odd.mem_bank[128],db_even.mem_bank[128],db_odd.mem_bank[129],db_even.mem_bank[129],db_odd.mem_bank[130],db_even.mem_bank[130],db_odd.mem_bank[131],db_even.mem_bank[131],db_odd.mem_bank[132],db_even.mem_bank[132],db_odd.mem_bank[133],db_even.mem_bank[133],db_odd.mem_bank[134],db_even.mem_bank[134],db_odd.mem_bank[135],db_even.mem_bank[135],db_odd.mem_bank[136],db_even.mem_bank[136],db_odd.mem_bank[137],db_even.mem_bank[137],db_odd.mem_bank[138],db_even.mem_bank[138],db_odd.mem_bank[139],db_even.mem_bank[139],db_odd.mem_bank[140],db_even.mem_bank[140],db_odd.mem_bank[141],db_even.mem_bank[141],db_odd.mem_bank[142],db_even.mem_bank[142],db_odd.mem_bank[143],db_even.mem_bank[143],db_odd.mem_bank[144],db_even.mem_bank[144],db_odd.mem_bank[145],db_even.mem_bank[145],db_odd.mem_bank[146],db_even.mem_bank[146],db_odd.mem_bank[147],db_even.mem_bank[147],db_odd.mem_bank[148],db_even.mem_bank[148],db_odd.mem_bank[149],db_even.mem_bank[149],db_odd.mem_bank[150],db_even.mem_bank[150],db_odd.mem_bank[151],db_even.mem_bank[151],db_odd.mem_bank[152],db_even.mem_bank[152],db_odd.mem_bank[153],db_even.mem_bank[153],db_odd.mem_bank[154],db_even.mem_bank[154],db_odd.mem_bank[155],db_even.mem_bank[155],db_odd.mem_bank[156],db_even.mem_bank[156],db_odd.mem_bank[157],db_even.mem_bank[157],db_odd.mem_bank[158],db_even.mem_bank[158],db_odd.mem_bank[159],db_even.mem_bank[159],db_odd.mem_bank[160],db_even.mem_bank[160],db_odd.mem_bank[161],db_even.mem_bank[161],db_odd.mem_bank[162],db_even.mem_bank[162],db_odd.mem_bank[163],db_even.mem_bank[163],db_odd.mem_bank[164],db_even.mem_bank[164],db_odd.mem_bank[165],db_even.mem_bank[165],db_odd.mem_bank[166],db_even.mem_bank[166],db_odd.mem_bank[167],db_even.mem_bank[167],db_odd.mem_bank[168],db_even.mem_bank[168],db_odd.mem_bank[169],db_even.mem_bank[169],db_odd.mem_bank[170],db_even.mem_bank[170],db_odd.mem_bank[171],db_even.mem_bank[171],db_odd.mem_bank[172],db_even.mem_bank[172],db_odd.mem_bank[173],db_even.mem_bank[173],db_odd.mem_bank[174],db_even.mem_bank[174],db_odd.mem_bank[175],db_even.mem_bank[175],db_odd.mem_bank[176],db_even.mem_bank[176],db_odd.mem_bank[177],db_even.mem_bank[177],db_odd.mem_bank[178],db_even.mem_bank[178],db_odd.mem_bank[179],db_even.mem_bank[179],db_odd.mem_bank[180],db_even.mem_bank[180],db_odd.mem_bank[181],db_even.mem_bank[181],db_odd.mem_bank[182],db_even.mem_bank[182],db_odd.mem_bank[183],db_even.mem_bank[183],db_odd.mem_bank[184],db_even.mem_bank[184],db_odd.mem_bank[185],db_even.mem_bank[185],db_odd.mem_bank[186],db_even.mem_bank[186],db_odd.mem_bank[187],db_even.mem_bank[187],db_odd.mem_bank[188],db_even.mem_bank[188],db_odd.mem_bank[189],db_even.mem_bank[189],db_odd.mem_bank[190],db_even.mem_bank[190],db_odd.mem_bank[191],db_even.mem_bank[191],db_odd.mem_bank[192],db_even.mem_bank[192],db_odd.mem_bank[193],db_even.mem_bank[193],db_odd.mem_bank[194],db_even.mem_bank[194],db_odd.mem_bank[195],db_even.mem_bank[195],db_odd.mem_bank[196],db_even.mem_bank[196],db_odd.mem_bank[197],db_even.mem_bank[197],db_odd.mem_bank[198],db_even.mem_bank[198],db_odd.mem_bank[199],db_even.mem_bank[199],db_odd.mem_bank[200],db_even.mem_bank[200],db_odd.mem_bank[201],db_even.mem_bank[201],db_odd.mem_bank[202],db_even.mem_bank[202],db_odd.mem_bank[203],db_even.mem_bank[203],db_odd.mem_bank[204],db_even.mem_bank[204],db_odd.mem_bank[205],db_even.mem_bank[205],db_odd.mem_bank[206],db_even.mem_bank[206],db_odd.mem_bank[207],db_even.mem_bank[207],db_odd.mem_bank[208],db_even.mem_bank[208],db_odd.mem_bank[209],db_even.mem_bank[209],db_odd.mem_bank[210],db_even.mem_bank[210],db_odd.mem_bank[211],db_even.mem_bank[211],db_odd.mem_bank[212],db_even.mem_bank[212],db_odd.mem_bank[213],db_even.mem_bank[213],db_odd.mem_bank[214],db_even.mem_bank[214],db_odd.mem_bank[215],db_even.mem_bank[215],db_odd.mem_bank[216],db_even.mem_bank[216],db_odd.mem_bank[217],db_even.mem_bank[217],db_odd.mem_bank[218],db_even.mem_bank[218],db_odd.mem_bank[219],db_even.mem_bank[219],db_odd.mem_bank[220],db_even.mem_bank[220],db_odd.mem_bank[221],db_even.mem_bank[221],db_odd.mem_bank[222],db_even.mem_bank[222],db_odd.mem_bank[223],db_even.mem_bank[223],db_odd.mem_bank[224],db_even.mem_bank[224],db_odd.mem_bank[225],db_even.mem_bank[225],db_odd.mem_bank[226],db_even.mem_bank[226],db_odd.mem_bank[227],db_even.mem_bank[227],db_odd.mem_bank[228],db_even.mem_bank[228],db_odd.mem_bank[229],db_even.mem_bank[229],db_odd.mem_bank[230],db_even.mem_bank[230],db_odd.mem_bank[231],db_even.mem_bank[231],db_odd.mem_bank[232],db_even.mem_bank[232],db_odd.mem_bank[233],db_even.mem_bank[233],db_odd.mem_bank[234],db_even.mem_bank[234],db_odd.mem_bank[235],db_even.mem_bank[235],db_odd.mem_bank[236],db_even.mem_bank[236],db_odd.mem_bank[237],db_even.mem_bank[237],db_odd.mem_bank[238],db_even.mem_bank[238],db_odd.mem_bank[239],db_even.mem_bank[239],db_odd.mem_bank[240],db_even.mem_bank[240],db_odd.mem_bank[241],db_even.mem_bank[241],db_odd.mem_bank[242],db_even.mem_bank[242],db_odd.mem_bank[243],db_even.mem_bank[243],db_odd.mem_bank[244],db_even.mem_bank[244],db_odd.mem_bank[245],db_even.mem_bank[245],db_odd.mem_bank[246],db_even.mem_bank[246],db_odd.mem_bank[247],db_even.mem_bank[247],db_odd.mem_bank[248],db_even.mem_bank[248],db_odd.mem_bank[249],db_even.mem_bank[249],db_odd.mem_bank[250],db_even.mem_bank[250],db_odd.mem_bank[251],db_even.mem_bank[251],db_odd.mem_bank[252],db_even.mem_bank[252],db_odd.mem_bank[253],db_even.mem_bank[253],db_odd.mem_bank[254],db_even.mem_bank[254],db_odd.mem_bank[255],db_even.mem_bank[255],db_odd.mem_bank[256],db_even.mem_bank[256],db_odd.mem_bank[257],db_even.mem_bank[257],db_odd.mem_bank[258],db_even.mem_bank[258],db_odd.mem_bank[259],db_even.mem_bank[259],db_odd.mem_bank[260],db_even.mem_bank[260],db_odd.mem_bank[261],db_even.mem_bank[261],db_odd.mem_bank[262],db_even.mem_bank[262],db_odd.mem_bank[263],db_even.mem_bank[263],db_odd.mem_bank[264],db_even.mem_bank[264],db_odd.mem_bank[265],db_even.mem_bank[265],db_odd.mem_bank[266],db_even.mem_bank[266],db_odd.mem_bank[267],db_even.mem_bank[267],db_odd.mem_bank[268],db_even.mem_bank[268],db_odd.mem_bank[269],db_even.mem_bank[269],db_odd.mem_bank[270],db_even.mem_bank[270],db_odd.mem_bank[271],db_even.mem_bank[271],db_odd.mem_bank[272],db_even.mem_bank[272],db_odd.mem_bank[273],db_even.mem_bank[273],db_odd.mem_bank[274],db_even.mem_bank[274],db_odd.mem_bank[275],db_even.mem_bank[275],db_odd.mem_bank[276],db_even.mem_bank[276],db_odd.mem_bank[277],db_even.mem_bank[277],db_odd.mem_bank[278],db_even.mem_bank[278],db_odd.mem_bank[279],db_even.mem_bank[279],db_odd.mem_bank[280],db_even.mem_bank[280],db_odd.mem_bank[281],db_even.mem_bank[281],db_odd.mem_bank[282],db_even.mem_bank[282],db_odd.mem_bank[283],db_even.mem_bank[283],db_odd.mem_bank[284],db_even.mem_bank[284],db_odd.mem_bank[285],db_even.mem_bank[285],db_odd.mem_bank[286],db_even.mem_bank[286],db_odd.mem_bank[287],db_even.mem_bank[287],db_odd.mem_bank[288],db_even.mem_bank[288],db_odd.mem_bank[289],db_even.mem_bank[289],db_odd.mem_bank[290],db_even.mem_bank[290],db_odd.mem_bank[291],db_even.mem_bank[291],db_odd.mem_bank[292],db_even.mem_bank[292],db_odd.mem_bank[293],db_even.mem_bank[293],db_odd.mem_bank[294],db_even.mem_bank[294],db_odd.mem_bank[295],db_even.mem_bank[295],db_odd.mem_bank[296],db_even.mem_bank[296],db_odd.mem_bank[297],db_even.mem_bank[297],db_odd.mem_bank[298],db_even.mem_bank[298],db_odd.mem_bank[299],db_even.mem_bank[299],db_odd.mem_bank[300],db_even.mem_bank[300],db_odd.mem_bank[301],db_even.mem_bank[301],db_odd.mem_bank[302],db_even.mem_bank[302],db_odd.mem_bank[303],db_even.mem_bank[303],db_odd.mem_bank[304],db_even.mem_bank[304],db_odd.mem_bank[305],db_even.mem_bank[305],db_odd.mem_bank[306],db_even.mem_bank[306],db_odd.mem_bank[307],db_even.mem_bank[307],db_odd.mem_bank[308],db_even.mem_bank[308],db_odd.mem_bank[309],db_even.mem_bank[309],db_odd.mem_bank[310],db_even.mem_bank[310],db_odd.mem_bank[311],db_even.mem_bank[311],db_odd.mem_bank[312],db_even.mem_bank[312],db_odd.mem_bank[313],db_even.mem_bank[313],db_odd.mem_bank[314],db_even.mem_bank[314],db_odd.mem_bank[315],db_even.mem_bank[315],db_odd.mem_bank[316],db_even.mem_bank[316],db_odd.mem_bank[317],db_even.mem_bank[317],db_odd.mem_bank[318],db_even.mem_bank[318],db_odd.mem_bank[319],db_even.mem_bank[319],db_odd.mem_bank[320],db_even.mem_bank[320],db_odd.mem_bank[321],db_even.mem_bank[321],db_odd.mem_bank[322],db_even.mem_bank[322],db_odd.mem_bank[323],db_even.mem_bank[323],db_odd.mem_bank[324],db_even.mem_bank[324],db_odd.mem_bank[325],db_even.mem_bank[325],db_odd.mem_bank[326],db_even.mem_bank[326],db_odd.mem_bank[327],db_even.mem_bank[327],db_odd.mem_bank[328],db_even.mem_bank[328],db_odd.mem_bank[329],db_even.mem_bank[329],db_odd.mem_bank[330],db_even.mem_bank[330],db_odd.mem_bank[331],db_even.mem_bank[331],db_odd.mem_bank[332],db_even.mem_bank[332],db_odd.mem_bank[333],db_even.mem_bank[333],db_odd.mem_bank[334],db_even.mem_bank[334],db_odd.mem_bank[335],db_even.mem_bank[335],db_odd.mem_bank[336],db_even.mem_bank[336],db_odd.mem_bank[337],db_even.mem_bank[337],db_odd.mem_bank[338],db_even.mem_bank[338],db_odd.mem_bank[339],db_even.mem_bank[339],db_odd.mem_bank[340],db_even.mem_bank[340],db_odd.mem_bank[341],db_even.mem_bank[341],db_odd.mem_bank[342],db_even.mem_bank[342],db_odd.mem_bank[343],db_even.mem_bank[343],db_odd.mem_bank[344],db_even.mem_bank[344],db_odd.mem_bank[345],db_even.mem_bank[345],db_odd.mem_bank[346],db_even.mem_bank[346],db_odd.mem_bank[347],db_even.mem_bank[347],db_odd.mem_bank[348],db_even.mem_bank[348],db_odd.mem_bank[349],db_even.mem_bank[349],db_odd.mem_bank[350],db_even.mem_bank[350],db_odd.mem_bank[351],db_even.mem_bank[351],db_odd.mem_bank[352],db_even.mem_bank[352],db_odd.mem_bank[353],db_even.mem_bank[353],db_odd.mem_bank[354],db_even.mem_bank[354],db_odd.mem_bank[355],db_even.mem_bank[355],db_odd.mem_bank[356],db_even.mem_bank[356],db_odd.mem_bank[357],db_even.mem_bank[357],db_odd.mem_bank[358],db_even.mem_bank[358],db_odd.mem_bank[359],db_even.mem_bank[359],db_odd.mem_bank[360],db_even.mem_bank[360],db_odd.mem_bank[361],db_even.mem_bank[361],db_odd.mem_bank[362],db_even.mem_bank[362],db_odd.mem_bank[363],db_even.mem_bank[363],db_odd.mem_bank[364],db_even.mem_bank[364],db_odd.mem_bank[365],db_even.mem_bank[365],db_odd.mem_bank[366],db_even.mem_bank[366],db_odd.mem_bank[367],db_even.mem_bank[367],db_odd.mem_bank[368],db_even.mem_bank[368],db_odd.mem_bank[369],db_even.mem_bank[369],db_odd.mem_bank[370],db_even.mem_bank[370],db_odd.mem_bank[371],db_even.mem_bank[371],db_odd.mem_bank[372],db_even.mem_bank[372],db_odd.mem_bank[373],db_even.mem_bank[373],db_odd.mem_bank[374],db_even.mem_bank[374],db_odd.mem_bank[375],db_even.mem_bank[375],db_odd.mem_bank[376],db_even.mem_bank[376],db_odd.mem_bank[377],db_even.mem_bank[377],db_odd.mem_bank[378],db_even.mem_bank[378],db_odd.mem_bank[379],db_even.mem_bank[379],db_odd.mem_bank[380],db_even.mem_bank[380],db_odd.mem_bank[381],db_even.mem_bank[381],db_odd.mem_bank[382],db_even.mem_bank[382],db_odd.mem_bank[383],db_even.mem_bank[383],db_odd.mem_bank[384],db_even.mem_bank[384],db_odd.mem_bank[385],db_even.mem_bank[385],db_odd.mem_bank[386],db_even.mem_bank[386],db_odd.mem_bank[387],db_even.mem_bank[387],db_odd.mem_bank[388],db_even.mem_bank[388],db_odd.mem_bank[389],db_even.mem_bank[389],db_odd.mem_bank[390],db_even.mem_bank[390],db_odd.mem_bank[391],db_even.mem_bank[391],db_odd.mem_bank[392],db_even.mem_bank[392],db_odd.mem_bank[393],db_even.mem_bank[393],db_odd.mem_bank[394],db_even.mem_bank[394],db_odd.mem_bank[395],db_even.mem_bank[395],db_odd.mem_bank[396],db_even.mem_bank[396],db_odd.mem_bank[397],db_even.mem_bank[397],db_odd.mem_bank[398],db_even.mem_bank[398],db_odd.mem_bank[399],db_even.mem_bank[399],db_odd.mem_bank[400],db_even.mem_bank[400],db_odd.mem_bank[401],db_even.mem_bank[401],db_odd.mem_bank[402],db_even.mem_bank[402],db_odd.mem_bank[403],db_even.mem_bank[403],db_odd.mem_bank[404],db_even.mem_bank[404],db_odd.mem_bank[405],db_even.mem_bank[405],db_odd.mem_bank[406],db_even.mem_bank[406],db_odd.mem_bank[407],db_even.mem_bank[407],db_odd.mem_bank[408],db_even.mem_bank[408],db_odd.mem_bank[409],db_even.mem_bank[409],db_odd.mem_bank[410],db_even.mem_bank[410],db_odd.mem_bank[411],db_even.mem_bank[411],db_odd.mem_bank[412],db_even.mem_bank[412],db_odd.mem_bank[413],db_even.mem_bank[413],db_odd.mem_bank[414],db_even.mem_bank[414],db_odd.mem_bank[415],db_even.mem_bank[415],db_odd.mem_bank[416],db_even.mem_bank[416],db_odd.mem_bank[417],db_even.mem_bank[417],db_odd.mem_bank[418],db_even.mem_bank[418],db_odd.mem_bank[419],db_even.mem_bank[419],db_odd.mem_bank[420],db_even.mem_bank[420],db_odd.mem_bank[421],db_even.mem_bank[421],db_odd.mem_bank[422],db_even.mem_bank[422],db_odd.mem_bank[423],db_even.mem_bank[423],db_odd.mem_bank[424],db_even.mem_bank[424],db_odd.mem_bank[425],db_even.mem_bank[425],db_odd.mem_bank[426],db_even.mem_bank[426],db_odd.mem_bank[427],db_even.mem_bank[427],db_odd.mem_bank[428],db_even.mem_bank[428],db_odd.mem_bank[429],db_even.mem_bank[429],db_odd.mem_bank[430],db_even.mem_bank[430],db_odd.mem_bank[431],db_even.mem_bank[431],db_odd.mem_bank[432],db_even.mem_bank[432],db_odd.mem_bank[433],db_even.mem_bank[433],db_odd.mem_bank[434],db_even.mem_bank[434],db_odd.mem_bank[435],db_even.mem_bank[435],db_odd.mem_bank[436],db_even.mem_bank[436],db_odd.mem_bank[437],db_even.mem_bank[437],db_odd.mem_bank[438],db_even.mem_bank[438],db_odd.mem_bank[439],db_even.mem_bank[439],db_odd.mem_bank[440],db_even.mem_bank[440],db_odd.mem_bank[441],db_even.mem_bank[441],db_odd.mem_bank[442],db_even.mem_bank[442],db_odd.mem_bank[443],db_even.mem_bank[443],db_odd.mem_bank[444],db_even.mem_bank[444],db_odd.mem_bank[445],db_even.mem_bank[445],db_odd.mem_bank[446],db_even.mem_bank[446],db_odd.mem_bank[447],db_even.mem_bank[447],db_odd.mem_bank[448],db_even.mem_bank[448],db_odd.mem_bank[449],db_even.mem_bank[449],db_odd.mem_bank[450],db_even.mem_bank[450],db_odd.mem_bank[451],db_even.mem_bank[451],db_odd.mem_bank[452],db_even.mem_bank[452],db_odd.mem_bank[453],db_even.mem_bank[453],db_odd.mem_bank[454],db_even.mem_bank[454],db_odd.mem_bank[455],db_even.mem_bank[455],db_odd.mem_bank[456],db_even.mem_bank[456],db_odd.mem_bank[457],db_even.mem_bank[457],db_odd.mem_bank[458],db_even.mem_bank[458],db_odd.mem_bank[459],db_even.mem_bank[459],db_odd.mem_bank[460],db_even.mem_bank[460],db_odd.mem_bank[461],db_even.mem_bank[461],db_odd.mem_bank[462],db_even.mem_bank[462],db_odd.mem_bank[463],db_even.mem_bank[463],db_odd.mem_bank[464],db_even.mem_bank[464],db_odd.mem_bank[465],db_even.mem_bank[465],db_odd.mem_bank[466],db_even.mem_bank[466],db_odd.mem_bank[467],db_even.mem_bank[467],db_odd.mem_bank[468],db_even.mem_bank[468],db_odd.mem_bank[469],db_even.mem_bank[469],db_odd.mem_bank[470],db_even.mem_bank[470],db_odd.mem_bank[471],db_even.mem_bank[471],db_odd.mem_bank[472],db_even.mem_bank[472],db_odd.mem_bank[473],db_even.mem_bank[473],db_odd.mem_bank[474],db_even.mem_bank[474],db_odd.mem_bank[475],db_even.mem_bank[475],db_odd.mem_bank[476],db_even.mem_bank[476],db_odd.mem_bank[477],db_even.mem_bank[477],db_odd.mem_bank[478],db_even.mem_bank[478],db_odd.mem_bank[479],db_even.mem_bank[479],db_odd.mem_bank[480],db_even.mem_bank[480],db_odd.mem_bank[481],db_even.mem_bank[481],db_odd.mem_bank[482],db_even.mem_bank[482],db_odd.mem_bank[483],db_even.mem_bank[483],db_odd.mem_bank[484],db_even.mem_bank[484],db_odd.mem_bank[485],db_even.mem_bank[485],db_odd.mem_bank[486],db_even.mem_bank[486],db_odd.mem_bank[487],db_even.mem_bank[487],db_odd.mem_bank[488],db_even.mem_bank[488],db_odd.mem_bank[489],db_even.mem_bank[489],db_odd.mem_bank[490],db_even.mem_bank[490],db_odd.mem_bank[491],db_even.mem_bank[491],db_odd.mem_bank[492],db_even.mem_bank[492],db_odd.mem_bank[493],db_even.mem_bank[493],db_odd.mem_bank[494],db_even.mem_bank[494],db_odd.mem_bank[495],db_even.mem_bank[495],db_odd.mem_bank[496],db_even.mem_bank[496],db_odd.mem_bank[497],db_even.mem_bank[497],db_odd.mem_bank[498],db_even.mem_bank[498],db_odd.mem_bank[499],db_even.mem_bank[499],db_odd.mem_bank[500],db_even.mem_bank[500],db_odd.mem_bank[501],db_even.mem_bank[501],db_odd.mem_bank[502],db_even.mem_bank[502],db_odd.mem_bank[503],db_even.mem_bank[503],db_odd.mem_bank[504],db_even.mem_bank[504],db_odd.mem_bank[505],db_even.mem_bank[505],db_odd.mem_bank[506],db_even.mem_bank[506],db_odd.mem_bank[507],db_even.mem_bank[507],db_odd.mem_bank[508],db_even.mem_bank[508],db_odd.mem_bank[509],db_even.mem_bank[509],db_odd.mem_bank[510],db_even.mem_bank[510],db_odd.mem_bank[511],db_even.mem_bank[511],db_odd.mem_bank[512],db_even.mem_bank[512],db_odd.mem_bank[513],db_even.mem_bank[513],db_odd.mem_bank[514],db_even.mem_bank[514],db_odd.mem_bank[515],db_even.mem_bank[515],db_odd.mem_bank[516],db_even.mem_bank[516],db_odd.mem_bank[517],db_even.mem_bank[517],db_odd.mem_bank[518],db_even.mem_bank[518],db_odd.mem_bank[519],db_even.mem_bank[519],db_odd.mem_bank[520],db_even.mem_bank[520],db_odd.mem_bank[521],db_even.mem_bank[521],db_odd.mem_bank[522],db_even.mem_bank[522],db_odd.mem_bank[523],db_even.mem_bank[523],db_odd.mem_bank[524],db_even.mem_bank[524],db_odd.mem_bank[525],db_even.mem_bank[525],db_odd.mem_bank[526],db_even.mem_bank[526],db_odd.mem_bank[527],db_even.mem_bank[527],db_odd.mem_bank[528],db_even.mem_bank[528],db_odd.mem_bank[529],db_even.mem_bank[529],db_odd.mem_bank[530],db_even.mem_bank[530],db_odd.mem_bank[531],db_even.mem_bank[531],db_odd.mem_bank[532],db_even.mem_bank[532],db_odd.mem_bank[533],db_even.mem_bank[533],db_odd.mem_bank[534],db_even.mem_bank[534],db_odd.mem_bank[535],db_even.mem_bank[535],db_odd.mem_bank[536],db_even.mem_bank[536],db_odd.mem_bank[537],db_even.mem_bank[537],db_odd.mem_bank[538],db_even.mem_bank[538],db_odd.mem_bank[539],db_even.mem_bank[539],db_odd.mem_bank[540],db_even.mem_bank[540],db_odd.mem_bank[541],db_even.mem_bank[541],db_odd.mem_bank[542],db_even.mem_bank[542],db_odd.mem_bank[543],db_even.mem_bank[543],db_odd.mem_bank[544],db_even.mem_bank[544],db_odd.mem_bank[545],db_even.mem_bank[545],db_odd.mem_bank[546],db_even.mem_bank[546],db_odd.mem_bank[547],db_even.mem_bank[547],db_odd.mem_bank[548],db_even.mem_bank[548],db_odd.mem_bank[549],db_even.mem_bank[549],db_odd.mem_bank[550],db_even.mem_bank[550],db_odd.mem_bank[551],db_even.mem_bank[551],db_odd.mem_bank[552],db_even.mem_bank[552],db_odd.mem_bank[553],db_even.mem_bank[553],db_odd.mem_bank[554],db_even.mem_bank[554],db_odd.mem_bank[555],db_even.mem_bank[555],db_odd.mem_bank[556],db_even.mem_bank[556],db_odd.mem_bank[557],db_even.mem_bank[557],db_odd.mem_bank[558],db_even.mem_bank[558],db_odd.mem_bank[559],db_even.mem_bank[559],db_odd.mem_bank[560],db_even.mem_bank[560],db_odd.mem_bank[561],db_even.mem_bank[561],db_odd.mem_bank[562],db_even.mem_bank[562],db_odd.mem_bank[563],db_even.mem_bank[563],db_odd.mem_bank[564],db_even.mem_bank[564],db_odd.mem_bank[565],db_even.mem_bank[565],db_odd.mem_bank[566],db_even.mem_bank[566],db_odd.mem_bank[567],db_even.mem_bank[567],db_odd.mem_bank[568],db_even.mem_bank[568],db_odd.mem_bank[569],db_even.mem_bank[569],db_odd.mem_bank[570],db_even.mem_bank[570],db_odd.mem_bank[571],db_even.mem_bank[571],db_odd.mem_bank[572],db_even.mem_bank[572],db_odd.mem_bank[573],db_even.mem_bank[573],db_odd.mem_bank[574],db_even.mem_bank[574],db_odd.mem_bank[575],db_even.mem_bank[575],db_odd.mem_bank[576],db_even.mem_bank[576],db_odd.mem_bank[577],db_even.mem_bank[577],db_odd.mem_bank[578],db_even.mem_bank[578],db_odd.mem_bank[579],db_even.mem_bank[579],db_odd.mem_bank[580],db_even.mem_bank[580],db_odd.mem_bank[581],db_even.mem_bank[581],db_odd.mem_bank[582],db_even.mem_bank[582],db_odd.mem_bank[583],db_even.mem_bank[583],db_odd.mem_bank[584],db_even.mem_bank[584],db_odd.mem_bank[585],db_even.mem_bank[585],db_odd.mem_bank[586],db_even.mem_bank[586],db_odd.mem_bank[587],db_even.mem_bank[587],db_odd.mem_bank[588],db_even.mem_bank[588],db_odd.mem_bank[589],db_even.mem_bank[589],db_odd.mem_bank[590],db_even.mem_bank[590],db_odd.mem_bank[591],db_even.mem_bank[591],db_odd.mem_bank[592],db_even.mem_bank[592],db_odd.mem_bank[593],db_even.mem_bank[593],db_odd.mem_bank[594],db_even.mem_bank[594],db_odd.mem_bank[595],db_even.mem_bank[595],db_odd.mem_bank[596],db_even.mem_bank[596],db_odd.mem_bank[597],db_even.mem_bank[597],db_odd.mem_bank[598],db_even.mem_bank[598],db_odd.mem_bank[599],db_even.mem_bank[599],db_odd.mem_bank[600],db_even.mem_bank[600],db_odd.mem_bank[601],db_even.mem_bank[601],db_odd.mem_bank[602],db_even.mem_bank[602],db_odd.mem_bank[603],db_even.mem_bank[603],db_odd.mem_bank[604],db_even.mem_bank[604],db_odd.mem_bank[605],db_even.mem_bank[605],db_odd.mem_bank[606],db_even.mem_bank[606],db_odd.mem_bank[607],db_even.mem_bank[607],db_odd.mem_bank[608],db_even.mem_bank[608],db_odd.mem_bank[609],db_even.mem_bank[609],db_odd.mem_bank[610],db_even.mem_bank[610],db_odd.mem_bank[611],db_even.mem_bank[611],db_odd.mem_bank[612],db_even.mem_bank[612],db_odd.mem_bank[613],db_even.mem_bank[613],db_odd.mem_bank[614],db_even.mem_bank[614],db_odd.mem_bank[615],db_even.mem_bank[615],db_odd.mem_bank[616],db_even.mem_bank[616],db_odd.mem_bank[617],db_even.mem_bank[617],db_odd.mem_bank[618],db_even.mem_bank[618],db_odd.mem_bank[619],db_even.mem_bank[619],db_odd.mem_bank[620],db_even.mem_bank[620],db_odd.mem_bank[621],db_even.mem_bank[621],db_odd.mem_bank[622],db_even.mem_bank[622],db_odd.mem_bank[623],db_even.mem_bank[623],db_odd.mem_bank[624],db_even.mem_bank[624],db_odd.mem_bank[625],db_even.mem_bank[625],db_odd.mem_bank[626],db_even.mem_bank[626],db_odd.mem_bank[627],db_even.mem_bank[627],db_odd.mem_bank[628],db_even.mem_bank[628],db_odd.mem_bank[629],db_even.mem_bank[629],db_odd.mem_bank[630],db_even.mem_bank[630],db_odd.mem_bank[631],db_even.mem_bank[631],db_odd.mem_bank[632],db_even.mem_bank[632],db_odd.mem_bank[633],db_even.mem_bank[633],db_odd.mem_bank[634],db_even.mem_bank[634],db_odd.mem_bank[635],db_even.mem_bank[635],db_odd.mem_bank[636],db_even.mem_bank[636],db_odd.mem_bank[637],db_even.mem_bank[637],db_odd.mem_bank[638],db_even.mem_bank[638],db_odd.mem_bank[639],db_even.mem_bank[639],db_odd.mem_bank[640],db_even.mem_bank[640],db_odd.mem_bank[641],db_even.mem_bank[641],db_odd.mem_bank[642],db_even.mem_bank[642],db_odd.mem_bank[643],db_even.mem_bank[643],db_odd.mem_bank[644],db_even.mem_bank[644],db_odd.mem_bank[645],db_even.mem_bank[645],db_odd.mem_bank[646],db_even.mem_bank[646],db_odd.mem_bank[647],db_even.mem_bank[647],db_odd.mem_bank[648],db_even.mem_bank[648],db_odd.mem_bank[649],db_even.mem_bank[649],db_odd.mem_bank[650],db_even.mem_bank[650],db_odd.mem_bank[651],db_even.mem_bank[651],db_odd.mem_bank[652],db_even.mem_bank[652],db_odd.mem_bank[653],db_even.mem_bank[653],db_odd.mem_bank[654],db_even.mem_bank[654],db_odd.mem_bank[655],db_even.mem_bank[655],db_odd.mem_bank[656],db_even.mem_bank[656],db_odd.mem_bank[657],db_even.mem_bank[657],db_odd.mem_bank[658],db_even.mem_bank[658],db_odd.mem_bank[659],db_even.mem_bank[659],db_odd.mem_bank[660],db_even.mem_bank[660],db_odd.mem_bank[661],db_even.mem_bank[661],db_odd.mem_bank[662],db_even.mem_bank[662],db_odd.mem_bank[663],db_even.mem_bank[663],db_odd.mem_bank[664],db_even.mem_bank[664],db_odd.mem_bank[665],db_even.mem_bank[665],db_odd.mem_bank[666],db_even.mem_bank[666],db_odd.mem_bank[667],db_even.mem_bank[667],db_odd.mem_bank[668],db_even.mem_bank[668],db_odd.mem_bank[669],db_even.mem_bank[669],db_odd.mem_bank[670],db_even.mem_bank[670],db_odd.mem_bank[671],db_even.mem_bank[671],db_odd.mem_bank[672],db_even.mem_bank[672],db_odd.mem_bank[673],db_even.mem_bank[673],db_odd.mem_bank[674],db_even.mem_bank[674],db_odd.mem_bank[675],db_even.mem_bank[675],db_odd.mem_bank[676],db_even.mem_bank[676],db_odd.mem_bank[677],db_even.mem_bank[677],db_odd.mem_bank[678],db_even.mem_bank[678],db_odd.mem_bank[679],db_even.mem_bank[679],db_odd.mem_bank[680],db_even.mem_bank[680],db_odd.mem_bank[681],db_even.mem_bank[681],db_odd.mem_bank[682],db_even.mem_bank[682],db_odd.mem_bank[683],db_even.mem_bank[683],db_odd.mem_bank[684],db_even.mem_bank[684],db_odd.mem_bank[685],db_even.mem_bank[685],db_odd.mem_bank[686],db_even.mem_bank[686],db_odd.mem_bank[687],db_even.mem_bank[687],db_odd.mem_bank[688],db_even.mem_bank[688],db_odd.mem_bank[689],db_even.mem_bank[689],db_odd.mem_bank[690],db_even.mem_bank[690],db_odd.mem_bank[691],db_even.mem_bank[691],db_odd.mem_bank[692],db_even.mem_bank[692],db_odd.mem_bank[693],db_even.mem_bank[693],db_odd.mem_bank[694],db_even.mem_bank[694],db_odd.mem_bank[695],db_even.mem_bank[695],db_odd.mem_bank[696],db_even.mem_bank[696],db_odd.mem_bank[697],db_even.mem_bank[697],db_odd.mem_bank[698],db_even.mem_bank[698],db_odd.mem_bank[699],db_even.mem_bank[699],db_odd.mem_bank[700],db_even.mem_bank[700],db_odd.mem_bank[701],db_even.mem_bank[701],db_odd.mem_bank[702],db_even.mem_bank[702],db_odd.mem_bank[703],db_even.mem_bank[703],db_odd.mem_bank[704],db_even.mem_bank[704],db_odd.mem_bank[705],db_even.mem_bank[705],db_odd.mem_bank[706],db_even.mem_bank[706],db_odd.mem_bank[707],db_even.mem_bank[707],db_odd.mem_bank[708],db_even.mem_bank[708],db_odd.mem_bank[709],db_even.mem_bank[709],db_odd.mem_bank[710],db_even.mem_bank[710],db_odd.mem_bank[711],db_even.mem_bank[711],db_odd.mem_bank[712],db_even.mem_bank[712],db_odd.mem_bank[713],db_even.mem_bank[713],db_odd.mem_bank[714],db_even.mem_bank[714],db_odd.mem_bank[715],db_even.mem_bank[715],db_odd.mem_bank[716],db_even.mem_bank[716],db_odd.mem_bank[717],db_even.mem_bank[717],db_odd.mem_bank[718],db_even.mem_bank[718],db_odd.mem_bank[719],db_even.mem_bank[719],db_odd.mem_bank[720],db_even.mem_bank[720],db_odd.mem_bank[721],db_even.mem_bank[721],db_odd.mem_bank[722],db_even.mem_bank[722],db_odd.mem_bank[723],db_even.mem_bank[723],db_odd.mem_bank[724],db_even.mem_bank[724],db_odd.mem_bank[725],db_even.mem_bank[725],db_odd.mem_bank[726],db_even.mem_bank[726],db_odd.mem_bank[727],db_even.mem_bank[727],db_odd.mem_bank[728],db_even.mem_bank[728],db_odd.mem_bank[729],db_even.mem_bank[729],db_odd.mem_bank[730],db_even.mem_bank[730],db_odd.mem_bank[731],db_even.mem_bank[731],db_odd.mem_bank[732],db_even.mem_bank[732],db_odd.mem_bank[733],db_even.mem_bank[733],db_odd.mem_bank[734],db_even.mem_bank[734],db_odd.mem_bank[735],db_even.mem_bank[735],db_odd.mem_bank[736],db_even.mem_bank[736],db_odd.mem_bank[737],db_even.mem_bank[737],db_odd.mem_bank[738],db_even.mem_bank[738],db_odd.mem_bank[739],db_even.mem_bank[739],db_odd.mem_bank[740],db_even.mem_bank[740],db_odd.mem_bank[741],db_even.mem_bank[741],db_odd.mem_bank[742],db_even.mem_bank[742],db_odd.mem_bank[743],db_even.mem_bank[743],db_odd.mem_bank[744],db_even.mem_bank[744],db_odd.mem_bank[745],db_even.mem_bank[745],db_odd.mem_bank[746],db_even.mem_bank[746],db_odd.mem_bank[747],db_even.mem_bank[747],db_odd.mem_bank[748],db_even.mem_bank[748],db_odd.mem_bank[749],db_even.mem_bank[749],db_odd.mem_bank[750],db_even.mem_bank[750],db_odd.mem_bank[751],db_even.mem_bank[751],db_odd.mem_bank[752],db_even.mem_bank[752],db_odd.mem_bank[753],db_even.mem_bank[753],db_odd.mem_bank[754],db_even.mem_bank[754],db_odd.mem_bank[755],db_even.mem_bank[755],db_odd.mem_bank[756],db_even.mem_bank[756],db_odd.mem_bank[757],db_even.mem_bank[757],db_odd.mem_bank[758],db_even.mem_bank[758],db_odd.mem_bank[759],db_even.mem_bank[759],db_odd.mem_bank[760],db_even.mem_bank[760],db_odd.mem_bank[761],db_even.mem_bank[761],db_odd.mem_bank[762],db_even.mem_bank[762],db_odd.mem_bank[763],db_even.mem_bank[763],db_odd.mem_bank[764],db_even.mem_bank[764],db_odd.mem_bank[765],db_even.mem_bank[765],db_odd.mem_bank[766],db_even.mem_bank[766],db_odd.mem_bank[767],db_even.mem_bank[767],db_odd.mem_bank[768],db_even.mem_bank[768],db_odd.mem_bank[769],db_even.mem_bank[769],db_odd.mem_bank[770],db_even.mem_bank[770],db_odd.mem_bank[771],db_even.mem_bank[771],db_odd.mem_bank[772],db_even.mem_bank[772],db_odd.mem_bank[773],db_even.mem_bank[773],db_odd.mem_bank[774],db_even.mem_bank[774],db_odd.mem_bank[775],db_even.mem_bank[775],db_odd.mem_bank[776],db_even.mem_bank[776],db_odd.mem_bank[777],db_even.mem_bank[777],db_odd.mem_bank[778],db_even.mem_bank[778],db_odd.mem_bank[779],db_even.mem_bank[779],db_odd.mem_bank[780],db_even.mem_bank[780],db_odd.mem_bank[781],db_even.mem_bank[781],db_odd.mem_bank[782],db_even.mem_bank[782],db_odd.mem_bank[783],db_even.mem_bank[783],db_odd.mem_bank[784],db_even.mem_bank[784],db_odd.mem_bank[785],db_even.mem_bank[785],db_odd.mem_bank[786],db_even.mem_bank[786],db_odd.mem_bank[787],db_even.mem_bank[787],db_odd.mem_bank[788],db_even.mem_bank[788],db_odd.mem_bank[789],db_even.mem_bank[789],db_odd.mem_bank[790],db_even.mem_bank[790],db_odd.mem_bank[791],db_even.mem_bank[791],db_odd.mem_bank[792],db_even.mem_bank[792],db_odd.mem_bank[793],db_even.mem_bank[793],db_odd.mem_bank[794],db_even.mem_bank[794],db_odd.mem_bank[795],db_even.mem_bank[795],db_odd.mem_bank[796],db_even.mem_bank[796],db_odd.mem_bank[797],db_even.mem_bank[797],db_odd.mem_bank[798],db_even.mem_bank[798],db_odd.mem_bank[799],db_even.mem_bank[799],db_odd.mem_bank[800],db_even.mem_bank[800],db_odd.mem_bank[801],db_even.mem_bank[801],db_odd.mem_bank[802],db_even.mem_bank[802],db_odd.mem_bank[803],db_even.mem_bank[803],db_odd.mem_bank[804],db_even.mem_bank[804],db_odd.mem_bank[805],db_even.mem_bank[805],db_odd.mem_bank[806],db_even.mem_bank[806],db_odd.mem_bank[807],db_even.mem_bank[807],db_odd.mem_bank[808],db_even.mem_bank[808],db_odd.mem_bank[809],db_even.mem_bank[809],db_odd.mem_bank[810],db_even.mem_bank[810],db_odd.mem_bank[811],db_even.mem_bank[811],db_odd.mem_bank[812],db_even.mem_bank[812],db_odd.mem_bank[813],db_even.mem_bank[813],db_odd.mem_bank[814],db_even.mem_bank[814],db_odd.mem_bank[815],db_even.mem_bank[815],db_odd.mem_bank[816],db_even.mem_bank[816],db_odd.mem_bank[817],db_even.mem_bank[817],db_odd.mem_bank[818],db_even.mem_bank[818],db_odd.mem_bank[819],db_even.mem_bank[819],db_odd.mem_bank[820],db_even.mem_bank[820],db_odd.mem_bank[821],db_even.mem_bank[821],db_odd.mem_bank[822],db_even.mem_bank[822],db_odd.mem_bank[823],db_even.mem_bank[823],db_odd.mem_bank[824],db_even.mem_bank[824],db_odd.mem_bank[825],db_even.mem_bank[825],db_odd.mem_bank[826],db_even.mem_bank[826],db_odd.mem_bank[827],db_even.mem_bank[827],db_odd.mem_bank[828],db_even.mem_bank[828],db_odd.mem_bank[829],db_even.mem_bank[829],db_odd.mem_bank[830],db_even.mem_bank[830],db_odd.mem_bank[831],db_even.mem_bank[831],db_odd.mem_bank[832],db_even.mem_bank[832],db_odd.mem_bank[833],db_even.mem_bank[833],db_odd.mem_bank[834],db_even.mem_bank[834],db_odd.mem_bank[835],db_even.mem_bank[835],db_odd.mem_bank[836],db_even.mem_bank[836],db_odd.mem_bank[837],db_even.mem_bank[837],db_odd.mem_bank[838],db_even.mem_bank[838],db_odd.mem_bank[839],db_even.mem_bank[839],db_odd.mem_bank[840],db_even.mem_bank[840],db_odd.mem_bank[841],db_even.mem_bank[841],db_odd.mem_bank[842],db_even.mem_bank[842],db_odd.mem_bank[843],db_even.mem_bank[843],db_odd.mem_bank[844],db_even.mem_bank[844],db_odd.mem_bank[845],db_even.mem_bank[845],db_odd.mem_bank[846],db_even.mem_bank[846],db_odd.mem_bank[847],db_even.mem_bank[847],db_odd.mem_bank[848],db_even.mem_bank[848],db_odd.mem_bank[849],db_even.mem_bank[849],db_odd.mem_bank[850],db_even.mem_bank[850],db_odd.mem_bank[851],db_even.mem_bank[851],db_odd.mem_bank[852],db_even.mem_bank[852],db_odd.mem_bank[853],db_even.mem_bank[853],db_odd.mem_bank[854],db_even.mem_bank[854],db_odd.mem_bank[855],db_even.mem_bank[855],db_odd.mem_bank[856],db_even.mem_bank[856],db_odd.mem_bank[857],db_even.mem_bank[857],db_odd.mem_bank[858],db_even.mem_bank[858],db_odd.mem_bank[859],db_even.mem_bank[859],db_odd.mem_bank[860],db_even.mem_bank[860],db_odd.mem_bank[861],db_even.mem_bank[861],db_odd.mem_bank[862],db_even.mem_bank[862],db_odd.mem_bank[863],db_even.mem_bank[863],db_odd.mem_bank[864],db_even.mem_bank[864],db_odd.mem_bank[865],db_even.mem_bank[865],db_odd.mem_bank[866],db_even.mem_bank[866],db_odd.mem_bank[867],db_even.mem_bank[867],db_odd.mem_bank[868],db_even.mem_bank[868],db_odd.mem_bank[869],db_even.mem_bank[869],db_odd.mem_bank[870],db_even.mem_bank[870],db_odd.mem_bank[871],db_even.mem_bank[871],db_odd.mem_bank[872],db_even.mem_bank[872],db_odd.mem_bank[873],db_even.mem_bank[873],db_odd.mem_bank[874],db_even.mem_bank[874],db_odd.mem_bank[875],db_even.mem_bank[875],db_odd.mem_bank[876],db_even.mem_bank[876],db_odd.mem_bank[877],db_even.mem_bank[877],db_odd.mem_bank[878],db_even.mem_bank[878],db_odd.mem_bank[879],db_even.mem_bank[879],db_odd.mem_bank[880],db_even.mem_bank[880],db_odd.mem_bank[881],db_even.mem_bank[881],db_odd.mem_bank[882],db_even.mem_bank[882],db_odd.mem_bank[883],db_even.mem_bank[883],db_odd.mem_bank[884],db_even.mem_bank[884],db_odd.mem_bank[885],db_even.mem_bank[885],db_odd.mem_bank[886],db_even.mem_bank[886],db_odd.mem_bank[887],db_even.mem_bank[887],db_odd.mem_bank[888],db_even.mem_bank[888],db_odd.mem_bank[889],db_even.mem_bank[889],db_odd.mem_bank[890],db_even.mem_bank[890],db_odd.mem_bank[891],db_even.mem_bank[891],db_odd.mem_bank[892],db_even.mem_bank[892],db_odd.mem_bank[893],db_even.mem_bank[893],db_odd.mem_bank[894],db_even.mem_bank[894],db_odd.mem_bank[895],db_even.mem_bank[895],db_odd.mem_bank[896],db_even.mem_bank[896],db_odd.mem_bank[897],db_even.mem_bank[897],db_odd.mem_bank[898],db_even.mem_bank[898],db_odd.mem_bank[899],db_even.mem_bank[899],db_odd.mem_bank[900],db_even.mem_bank[900],db_odd.mem_bank[901],db_even.mem_bank[901],db_odd.mem_bank[902],db_even.mem_bank[902],db_odd.mem_bank[903],db_even.mem_bank[903],db_odd.mem_bank[904],db_even.mem_bank[904],db_odd.mem_bank[905],db_even.mem_bank[905],db_odd.mem_bank[906],db_even.mem_bank[906],db_odd.mem_bank[907],db_even.mem_bank[907],db_odd.mem_bank[908],db_even.mem_bank[908],db_odd.mem_bank[909],db_even.mem_bank[909],db_odd.mem_bank[910],db_even.mem_bank[910],db_odd.mem_bank[911],db_even.mem_bank[911],db_odd.mem_bank[912],db_even.mem_bank[912],db_odd.mem_bank[913],db_even.mem_bank[913],db_odd.mem_bank[914],db_even.mem_bank[914],db_odd.mem_bank[915],db_even.mem_bank[915],db_odd.mem_bank[916],db_even.mem_bank[916],db_odd.mem_bank[917],db_even.mem_bank[917],db_odd.mem_bank[918],db_even.mem_bank[918],db_odd.mem_bank[919],db_even.mem_bank[919],db_odd.mem_bank[920],db_even.mem_bank[920],db_odd.mem_bank[921],db_even.mem_bank[921],db_odd.mem_bank[922],db_even.mem_bank[922],db_odd.mem_bank[923],db_even.mem_bank[923],db_odd.mem_bank[924],db_even.mem_bank[924],db_odd.mem_bank[925],db_even.mem_bank[925],db_odd.mem_bank[926],db_even.mem_bank[926],db_odd.mem_bank[927],db_even.mem_bank[927],db_odd.mem_bank[928],db_even.mem_bank[928],db_odd.mem_bank[929],db_even.mem_bank[929],db_odd.mem_bank[930],db_even.mem_bank[930],db_odd.mem_bank[931],db_even.mem_bank[931],db_odd.mem_bank[932],db_even.mem_bank[932],db_odd.mem_bank[933],db_even.mem_bank[933],db_odd.mem_bank[934],db_even.mem_bank[934],db_odd.mem_bank[935],db_even.mem_bank[935],db_odd.mem_bank[936],db_even.mem_bank[936],db_odd.mem_bank[937],db_even.mem_bank[937],db_odd.mem_bank[938],db_even.mem_bank[938],db_odd.mem_bank[939],db_even.mem_bank[939],db_odd.mem_bank[940],db_even.mem_bank[940],db_odd.mem_bank[941],db_even.mem_bank[941],db_odd.mem_bank[942],db_even.mem_bank[942],db_odd.mem_bank[943],db_even.mem_bank[943],db_odd.mem_bank[944],db_even.mem_bank[944],db_odd.mem_bank[945],db_even.mem_bank[945],db_odd.mem_bank[946],db_even.mem_bank[946],db_odd.mem_bank[947],db_even.mem_bank[947],db_odd.mem_bank[948],db_even.mem_bank[948],db_odd.mem_bank[949],db_even.mem_bank[949],db_odd.mem_bank[950],db_even.mem_bank[950],db_odd.mem_bank[951],db_even.mem_bank[951],db_odd.mem_bank[952],db_even.mem_bank[952],db_odd.mem_bank[953],db_even.mem_bank[953],db_odd.mem_bank[954],db_even.mem_bank[954],db_odd.mem_bank[955],db_even.mem_bank[955],db_odd.mem_bank[956],db_even.mem_bank[956],db_odd.mem_bank[957],db_even.mem_bank[957],db_odd.mem_bank[958],db_even.mem_bank[958],db_odd.mem_bank[959],db_even.mem_bank[959],db_odd.mem_bank[960],db_even.mem_bank[960],db_odd.mem_bank[961],db_even.mem_bank[961],db_odd.mem_bank[962],db_even.mem_bank[962],db_odd.mem_bank[963],db_even.mem_bank[963],db_odd.mem_bank[964],db_even.mem_bank[964],db_odd.mem_bank[965],db_even.mem_bank[965],db_odd.mem_bank[966],db_even.mem_bank[966],db_odd.mem_bank[967],db_even.mem_bank[967],db_odd.mem_bank[968],db_even.mem_bank[968],db_odd.mem_bank[969],db_even.mem_bank[969],db_odd.mem_bank[970],db_even.mem_bank[970],db_odd.mem_bank[971],db_even.mem_bank[971],db_odd.mem_bank[972],db_even.mem_bank[972],db_odd.mem_bank[973],db_even.mem_bank[973],db_odd.mem_bank[974],db_even.mem_bank[974],db_odd.mem_bank[975],db_even.mem_bank[975],db_odd.mem_bank[976],db_even.mem_bank[976],db_odd.mem_bank[977],db_even.mem_bank[977],db_odd.mem_bank[978],db_even.mem_bank[978],db_odd.mem_bank[979],db_even.mem_bank[979],db_odd.mem_bank[980],db_even.mem_bank[980],db_odd.mem_bank[981],db_even.mem_bank[981],db_odd.mem_bank[982],db_even.mem_bank[982],db_odd.mem_bank[983],db_even.mem_bank[983],db_odd.mem_bank[984],db_even.mem_bank[984],db_odd.mem_bank[985],db_even.mem_bank[985],db_odd.mem_bank[986],db_even.mem_bank[986],db_odd.mem_bank[987],db_even.mem_bank[987],db_odd.mem_bank[988],db_even.mem_bank[988],db_odd.mem_bank[989],db_even.mem_bank[989],db_odd.mem_bank[990],db_even.mem_bank[990],db_odd.mem_bank[991],db_even.mem_bank[991],db_odd.mem_bank[992],db_even.mem_bank[992],db_odd.mem_bank[993],db_even.mem_bank[993],db_odd.mem_bank[994],db_even.mem_bank[994],db_odd.mem_bank[995],db_even.mem_bank[995],db_odd.mem_bank[996],db_even.mem_bank[996],db_odd.mem_bank[997],db_even.mem_bank[997],db_odd.mem_bank[998],db_even.mem_bank[998],db_odd.mem_bank[999],db_even.mem_bank[999],db_odd.mem_bank[1000],db_even.mem_bank[1000],db_odd.mem_bank[1001],db_even.mem_bank[1001],db_odd.mem_bank[1002],db_even.mem_bank[1002],db_odd.mem_bank[1003],db_even.mem_bank[1003],db_odd.mem_bank[1004],db_even.mem_bank[1004],db_odd.mem_bank[1005],db_even.mem_bank[1005],db_odd.mem_bank[1006],db_even.mem_bank[1006],db_odd.mem_bank[1007],db_even.mem_bank[1007],db_odd.mem_bank[1008],db_even.mem_bank[1008],db_odd.mem_bank[1009],db_even.mem_bank[1009],db_odd.mem_bank[1010],db_even.mem_bank[1010],db_odd.mem_bank[1011],db_even.mem_bank[1011],db_odd.mem_bank[1012],db_even.mem_bank[1012],db_odd.mem_bank[1013],db_even.mem_bank[1013],db_odd.mem_bank[1014],db_even.mem_bank[1014],db_odd.mem_bank[1015],db_even.mem_bank[1015],db_odd.mem_bank[1016],db_even.mem_bank[1016],db_odd.mem_bank[1017],db_even.mem_bank[1017],db_odd.mem_bank[1018],db_even.mem_bank[1018],db_odd.mem_bank[1019],db_even.mem_bank[1019],db_odd.mem_bank[1020],db_even.mem_bank[1020],db_odd.mem_bank[1021],db_even.mem_bank[1021],db_odd.mem_bank[1022],db_even.mem_bank[1022],db_odd.mem_bank[1023],db_even.mem_bank[1023],db_odd.mem_bank[1024],db_even.mem_bank[1024],db_odd.mem_bank[1025],db_even.mem_bank[1025],db_odd.mem_bank[1026],db_even.mem_bank[1026],db_odd.mem_bank[1027],db_even.mem_bank[1027],db_odd.mem_bank[1028],db_even.mem_bank[1028],db_odd.mem_bank[1029],db_even.mem_bank[1029],db_odd.mem_bank[1030],db_even.mem_bank[1030],db_odd.mem_bank[1031],db_even.mem_bank[1031],db_odd.mem_bank[1032],db_even.mem_bank[1032],db_odd.mem_bank[1033],db_even.mem_bank[1033],db_odd.mem_bank[1034],db_even.mem_bank[1034],db_odd.mem_bank[1035],db_even.mem_bank[1035],db_odd.mem_bank[1036],db_even.mem_bank[1036],db_odd.mem_bank[1037],db_even.mem_bank[1037],db_odd.mem_bank[1038],db_even.mem_bank[1038],db_odd.mem_bank[1039],db_even.mem_bank[1039],db_odd.mem_bank[1040],db_even.mem_bank[1040],db_odd.mem_bank[1041],db_even.mem_bank[1041],db_odd.mem_bank[1042],db_even.mem_bank[1042],db_odd.mem_bank[1043],db_even.mem_bank[1043],db_odd.mem_bank[1044],db_even.mem_bank[1044],db_odd.mem_bank[1045],db_even.mem_bank[1045],db_odd.mem_bank[1046],db_even.mem_bank[1046],db_odd.mem_bank[1047],db_even.mem_bank[1047],db_odd.mem_bank[1048],db_even.mem_bank[1048],db_odd.mem_bank[1049],db_even.mem_bank[1049],db_odd.mem_bank[1050],db_even.mem_bank[1050],db_odd.mem_bank[1051],db_even.mem_bank[1051],db_odd.mem_bank[1052],db_even.mem_bank[1052],db_odd.mem_bank[1053],db_even.mem_bank[1053],db_odd.mem_bank[1054],db_even.mem_bank[1054],db_odd.mem_bank[1055],db_even.mem_bank[1055],db_odd.mem_bank[1056],db_even.mem_bank[1056],db_odd.mem_bank[1057],db_even.mem_bank[1057],db_odd.mem_bank[1058],db_even.mem_bank[1058],db_odd.mem_bank[1059],db_even.mem_bank[1059],db_odd.mem_bank[1060],db_even.mem_bank[1060],db_odd.mem_bank[1061],db_even.mem_bank[1061],db_odd.mem_bank[1062],db_even.mem_bank[1062],db_odd.mem_bank[1063],db_even.mem_bank[1063],db_odd.mem_bank[1064],db_even.mem_bank[1064],db_odd.mem_bank[1065],db_even.mem_bank[1065],db_odd.mem_bank[1066],db_even.mem_bank[1066],db_odd.mem_bank[1067],db_even.mem_bank[1067],db_odd.mem_bank[1068],db_even.mem_bank[1068],db_odd.mem_bank[1069],db_even.mem_bank[1069],db_odd.mem_bank[1070],db_even.mem_bank[1070],db_odd.mem_bank[1071],db_even.mem_bank[1071],db_odd.mem_bank[1072],db_even.mem_bank[1072],db_odd.mem_bank[1073],db_even.mem_bank[1073],db_odd.mem_bank[1074],db_even.mem_bank[1074],db_odd.mem_bank[1075],db_even.mem_bank[1075],db_odd.mem_bank[1076],db_even.mem_bank[1076],db_odd.mem_bank[1077],db_even.mem_bank[1077],db_odd.mem_bank[1078],db_even.mem_bank[1078],db_odd.mem_bank[1079],db_even.mem_bank[1079],db_odd.mem_bank[1080],db_even.mem_bank[1080],db_odd.mem_bank[1081],db_even.mem_bank[1081],db_odd.mem_bank[1082],db_even.mem_bank[1082],db_odd.mem_bank[1083],db_even.mem_bank[1083],db_odd.mem_bank[1084],db_even.mem_bank[1084],db_odd.mem_bank[1085],db_even.mem_bank[1085],db_odd.mem_bank[1086],db_even.mem_bank[1086],db_odd.mem_bank[1087],db_even.mem_bank[1087],db_odd.mem_bank[1088],db_even.mem_bank[1088],db_odd.mem_bank[1089],db_even.mem_bank[1089],db_odd.mem_bank[1090],db_even.mem_bank[1090],db_odd.mem_bank[1091],db_even.mem_bank[1091],db_odd.mem_bank[1092],db_even.mem_bank[1092],db_odd.mem_bank[1093],db_even.mem_bank[1093],db_odd.mem_bank[1094],db_even.mem_bank[1094],db_odd.mem_bank[1095],db_even.mem_bank[1095],db_odd.mem_bank[1096],db_even.mem_bank[1096],db_odd.mem_bank[1097],db_even.mem_bank[1097],db_odd.mem_bank[1098],db_even.mem_bank[1098],db_odd.mem_bank[1099],db_even.mem_bank[1099],db_odd.mem_bank[1100],db_even.mem_bank[1100],db_odd.mem_bank[1101],db_even.mem_bank[1101],db_odd.mem_bank[1102],db_even.mem_bank[1102],db_odd.mem_bank[1103],db_even.mem_bank[1103],db_odd.mem_bank[1104],db_even.mem_bank[1104],db_odd.mem_bank[1105],db_even.mem_bank[1105],db_odd.mem_bank[1106],db_even.mem_bank[1106],db_odd.mem_bank[1107],db_even.mem_bank[1107],db_odd.mem_bank[1108],db_even.mem_bank[1108],db_odd.mem_bank[1109],db_even.mem_bank[1109],db_odd.mem_bank[1110],db_even.mem_bank[1110],db_odd.mem_bank[1111],db_even.mem_bank[1111],db_odd.mem_bank[1112],db_even.mem_bank[1112],db_odd.mem_bank[1113],db_even.mem_bank[1113],db_odd.mem_bank[1114],db_even.mem_bank[1114],db_odd.mem_bank[1115],db_even.mem_bank[1115],db_odd.mem_bank[1116],db_even.mem_bank[1116],db_odd.mem_bank[1117],db_even.mem_bank[1117],db_odd.mem_bank[1118],db_even.mem_bank[1118],db_odd.mem_bank[1119],db_even.mem_bank[1119],db_odd.mem_bank[1120],db_even.mem_bank[1120],db_odd.mem_bank[1121],db_even.mem_bank[1121],db_odd.mem_bank[1122],db_even.mem_bank[1122],db_odd.mem_bank[1123],db_even.mem_bank[1123],db_odd.mem_bank[1124],db_even.mem_bank[1124],db_odd.mem_bank[1125],db_even.mem_bank[1125],db_odd.mem_bank[1126],db_even.mem_bank[1126],db_odd.mem_bank[1127],db_even.mem_bank[1127],db_odd.mem_bank[1128],db_even.mem_bank[1128],db_odd.mem_bank[1129],db_even.mem_bank[1129],db_odd.mem_bank[1130],db_even.mem_bank[1130],db_odd.mem_bank[1131],db_even.mem_bank[1131],db_odd.mem_bank[1132],db_even.mem_bank[1132],db_odd.mem_bank[1133],db_even.mem_bank[1133],db_odd.mem_bank[1134],db_even.mem_bank[1134],db_odd.mem_bank[1135],db_even.mem_bank[1135],db_odd.mem_bank[1136],db_even.mem_bank[1136],db_odd.mem_bank[1137],db_even.mem_bank[1137],db_odd.mem_bank[1138],db_even.mem_bank[1138],db_odd.mem_bank[1139],db_even.mem_bank[1139],db_odd.mem_bank[1140],db_even.mem_bank[1140],db_odd.mem_bank[1141],db_even.mem_bank[1141],db_odd.mem_bank[1142],db_even.mem_bank[1142],db_odd.mem_bank[1143],db_even.mem_bank[1143],db_odd.mem_bank[1144],db_even.mem_bank[1144],db_odd.mem_bank[1145],db_even.mem_bank[1145],db_odd.mem_bank[1146],db_even.mem_bank[1146],db_odd.mem_bank[1147],db_even.mem_bank[1147],db_odd.mem_bank[1148],db_even.mem_bank[1148],db_odd.mem_bank[1149],db_even.mem_bank[1149],db_odd.mem_bank[1150],db_even.mem_bank[1150],db_odd.mem_bank[1151],db_even.mem_bank[1151],db_odd.mem_bank[1152],db_even.mem_bank[1152],db_odd.mem_bank[1153],db_even.mem_bank[1153],db_odd.mem_bank[1154],db_even.mem_bank[1154],db_odd.mem_bank[1155],db_even.mem_bank[1155],db_odd.mem_bank[1156],db_even.mem_bank[1156],db_odd.mem_bank[1157],db_even.mem_bank[1157],db_odd.mem_bank[1158],db_even.mem_bank[1158],db_odd.mem_bank[1159],db_even.mem_bank[1159],db_odd.mem_bank[1160],db_even.mem_bank[1160],db_odd.mem_bank[1161],db_even.mem_bank[1161],db_odd.mem_bank[1162],db_even.mem_bank[1162],db_odd.mem_bank[1163],db_even.mem_bank[1163],db_odd.mem_bank[1164],db_even.mem_bank[1164],db_odd.mem_bank[1165],db_even.mem_bank[1165],db_odd.mem_bank[1166],db_even.mem_bank[1166],db_odd.mem_bank[1167],db_even.mem_bank[1167],db_odd.mem_bank[1168],db_even.mem_bank[1168],db_odd.mem_bank[1169],db_even.mem_bank[1169],db_odd.mem_bank[1170],db_even.mem_bank[1170],db_odd.mem_bank[1171],db_even.mem_bank[1171],db_odd.mem_bank[1172],db_even.mem_bank[1172],db_odd.mem_bank[1173],db_even.mem_bank[1173],db_odd.mem_bank[1174],db_even.mem_bank[1174],db_odd.mem_bank[1175],db_even.mem_bank[1175],db_odd.mem_bank[1176],db_even.mem_bank[1176],db_odd.mem_bank[1177],db_even.mem_bank[1177],db_odd.mem_bank[1178],db_even.mem_bank[1178],db_odd.mem_bank[1179],db_even.mem_bank[1179],db_odd.mem_bank[1180],db_even.mem_bank[1180],db_odd.mem_bank[1181],db_even.mem_bank[1181],db_odd.mem_bank[1182],db_even.mem_bank[1182],db_odd.mem_bank[1183],db_even.mem_bank[1183],db_odd.mem_bank[1184],db_even.mem_bank[1184],db_odd.mem_bank[1185],db_even.mem_bank[1185],db_odd.mem_bank[1186],db_even.mem_bank[1186],db_odd.mem_bank[1187],db_even.mem_bank[1187],db_odd.mem_bank[1188],db_even.mem_bank[1188],db_odd.mem_bank[1189],db_even.mem_bank[1189],db_odd.mem_bank[1190],db_even.mem_bank[1190],db_odd.mem_bank[1191],db_even.mem_bank[1191],db_odd.mem_bank[1192],db_even.mem_bank[1192],db_odd.mem_bank[1193],db_even.mem_bank[1193],db_odd.mem_bank[1194],db_even.mem_bank[1194],db_odd.mem_bank[1195],db_even.mem_bank[1195],db_odd.mem_bank[1196],db_even.mem_bank[1196],db_odd.mem_bank[1197],db_even.mem_bank[1197],db_odd.mem_bank[1198],db_even.mem_bank[1198],db_odd.mem_bank[1199],db_even.mem_bank[1199],db_odd.mem_bank[1200],db_even.mem_bank[1200],db_odd.mem_bank[1201],db_even.mem_bank[1201],db_odd.mem_bank[1202],db_even.mem_bank[1202],db_odd.mem_bank[1203],db_even.mem_bank[1203],db_odd.mem_bank[1204],db_even.mem_bank[1204],db_odd.mem_bank[1205],db_even.mem_bank[1205],db_odd.mem_bank[1206],db_even.mem_bank[1206],db_odd.mem_bank[1207],db_even.mem_bank[1207],db_odd.mem_bank[1208],db_even.mem_bank[1208],db_odd.mem_bank[1209],db_even.mem_bank[1209],db_odd.mem_bank[1210],db_even.mem_bank[1210],db_odd.mem_bank[1211],db_even.mem_bank[1211],db_odd.mem_bank[1212],db_even.mem_bank[1212],db_odd.mem_bank[1213],db_even.mem_bank[1213],db_odd.mem_bank[1214],db_even.mem_bank[1214],db_odd.mem_bank[1215],db_even.mem_bank[1215],db_odd.mem_bank[1216],db_even.mem_bank[1216],db_odd.mem_bank[1217],db_even.mem_bank[1217],db_odd.mem_bank[1218],db_even.mem_bank[1218],db_odd.mem_bank[1219],db_even.mem_bank[1219],db_odd.mem_bank[1220],db_even.mem_bank[1220],db_odd.mem_bank[1221],db_even.mem_bank[1221],db_odd.mem_bank[1222],db_even.mem_bank[1222],db_odd.mem_bank[1223],db_even.mem_bank[1223],db_odd.mem_bank[1224],db_even.mem_bank[1224],db_odd.mem_bank[1225],db_even.mem_bank[1225],db_odd.mem_bank[1226],db_even.mem_bank[1226],db_odd.mem_bank[1227],db_even.mem_bank[1227],db_odd.mem_bank[1228],db_even.mem_bank[1228],db_odd.mem_bank[1229],db_even.mem_bank[1229],db_odd.mem_bank[1230],db_even.mem_bank[1230],db_odd.mem_bank[1231],db_even.mem_bank[1231],db_odd.mem_bank[1232],db_even.mem_bank[1232],db_odd.mem_bank[1233],db_even.mem_bank[1233],db_odd.mem_bank[1234],db_even.mem_bank[1234],db_odd.mem_bank[1235],db_even.mem_bank[1235],db_odd.mem_bank[1236],db_even.mem_bank[1236],db_odd.mem_bank[1237],db_even.mem_bank[1237],db_odd.mem_bank[1238],db_even.mem_bank[1238],db_odd.mem_bank[1239],db_even.mem_bank[1239],db_odd.mem_bank[1240],db_even.mem_bank[1240],db_odd.mem_bank[1241],db_even.mem_bank[1241],db_odd.mem_bank[1242],db_even.mem_bank[1242],db_odd.mem_bank[1243],db_even.mem_bank[1243],db_odd.mem_bank[1244],db_even.mem_bank[1244],db_odd.mem_bank[1245],db_even.mem_bank[1245],db_odd.mem_bank[1246],db_even.mem_bank[1246],db_odd.mem_bank[1247],db_even.mem_bank[1247],db_odd.mem_bank[1248],db_even.mem_bank[1248],db_odd.mem_bank[1249],db_even.mem_bank[1249],db_odd.mem_bank[1250],db_even.mem_bank[1250],db_odd.mem_bank[1251],db_even.mem_bank[1251],db_odd.mem_bank[1252],db_even.mem_bank[1252],db_odd.mem_bank[1253],db_even.mem_bank[1253],db_odd.mem_bank[1254],db_even.mem_bank[1254],db_odd.mem_bank[1255],db_even.mem_bank[1255],db_odd.mem_bank[1256],db_even.mem_bank[1256],db_odd.mem_bank[1257],db_even.mem_bank[1257],db_odd.mem_bank[1258],db_even.mem_bank[1258],db_odd.mem_bank[1259],db_even.mem_bank[1259],db_odd.mem_bank[1260],db_even.mem_bank[1260],db_odd.mem_bank[1261],db_even.mem_bank[1261],db_odd.mem_bank[1262],db_even.mem_bank[1262],db_odd.mem_bank[1263],db_even.mem_bank[1263],db_odd.mem_bank[1264],db_even.mem_bank[1264],db_odd.mem_bank[1265],db_even.mem_bank[1265],db_odd.mem_bank[1266],db_even.mem_bank[1266],db_odd.mem_bank[1267],db_even.mem_bank[1267],db_odd.mem_bank[1268],db_even.mem_bank[1268],db_odd.mem_bank[1269],db_even.mem_bank[1269],db_odd.mem_bank[1270],db_even.mem_bank[1270],db_odd.mem_bank[1271],db_even.mem_bank[1271],db_odd.mem_bank[1272],db_even.mem_bank[1272],db_odd.mem_bank[1273],db_even.mem_bank[1273],db_odd.mem_bank[1274],db_even.mem_bank[1274],db_odd.mem_bank[1275],db_even.mem_bank[1275],db_odd.mem_bank[1276],db_even.mem_bank[1276],db_odd.mem_bank[1277],db_even.mem_bank[1277],db_odd.mem_bank[1278],db_even.mem_bank[1278],db_odd.mem_bank[1279],db_even.mem_bank[1279],db_odd.mem_bank[1280],db_even.mem_bank[1280],db_odd.mem_bank[1281],db_even.mem_bank[1281],db_odd.mem_bank[1282],db_even.mem_bank[1282],db_odd.mem_bank[1283],db_even.mem_bank[1283],db_odd.mem_bank[1284],db_even.mem_bank[1284],db_odd.mem_bank[1285],db_even.mem_bank[1285],db_odd.mem_bank[1286],db_even.mem_bank[1286],db_odd.mem_bank[1287],db_even.mem_bank[1287],db_odd.mem_bank[1288],db_even.mem_bank[1288],db_odd.mem_bank[1289],db_even.mem_bank[1289],db_odd.mem_bank[1290],db_even.mem_bank[1290],db_odd.mem_bank[1291],db_even.mem_bank[1291],db_odd.mem_bank[1292],db_even.mem_bank[1292],db_odd.mem_bank[1293],db_even.mem_bank[1293],db_odd.mem_bank[1294],db_even.mem_bank[1294],db_odd.mem_bank[1295],db_even.mem_bank[1295],db_odd.mem_bank[1296],db_even.mem_bank[1296],db_odd.mem_bank[1297],db_even.mem_bank[1297],db_odd.mem_bank[1298],db_even.mem_bank[1298],db_odd.mem_bank[1299],db_even.mem_bank[1299],db_odd.mem_bank[1300],db_even.mem_bank[1300],db_odd.mem_bank[1301],db_even.mem_bank[1301],db_odd.mem_bank[1302],db_even.mem_bank[1302],db_odd.mem_bank[1303],db_even.mem_bank[1303],db_odd.mem_bank[1304],db_even.mem_bank[1304],db_odd.mem_bank[1305],db_even.mem_bank[1305],db_odd.mem_bank[1306],db_even.mem_bank[1306],db_odd.mem_bank[1307],db_even.mem_bank[1307],db_odd.mem_bank[1308],db_even.mem_bank[1308],db_odd.mem_bank[1309],db_even.mem_bank[1309],db_odd.mem_bank[1310],db_even.mem_bank[1310],db_odd.mem_bank[1311],db_even.mem_bank[1311],db_odd.mem_bank[1312],db_even.mem_bank[1312],db_odd.mem_bank[1313],db_even.mem_bank[1313],db_odd.mem_bank[1314],db_even.mem_bank[1314],db_odd.mem_bank[1315],db_even.mem_bank[1315],db_odd.mem_bank[1316],db_even.mem_bank[1316],db_odd.mem_bank[1317],db_even.mem_bank[1317],db_odd.mem_bank[1318],db_even.mem_bank[1318],db_odd.mem_bank[1319],db_even.mem_bank[1319],db_odd.mem_bank[1320],db_even.mem_bank[1320],db_odd.mem_bank[1321],db_even.mem_bank[1321],db_odd.mem_bank[1322],db_even.mem_bank[1322],db_odd.mem_bank[1323],db_even.mem_bank[1323],db_odd.mem_bank[1324],db_even.mem_bank[1324],db_odd.mem_bank[1325],db_even.mem_bank[1325],db_odd.mem_bank[1326],db_even.mem_bank[1326],db_odd.mem_bank[1327],db_even.mem_bank[1327],db_odd.mem_bank[1328],db_even.mem_bank[1328],db_odd.mem_bank[1329],db_even.mem_bank[1329],db_odd.mem_bank[1330],db_even.mem_bank[1330],db_odd.mem_bank[1331],db_even.mem_bank[1331],db_odd.mem_bank[1332],db_even.mem_bank[1332],db_odd.mem_bank[1333],db_even.mem_bank[1333],db_odd.mem_bank[1334],db_even.mem_bank[1334],db_odd.mem_bank[1335],db_even.mem_bank[1335],db_odd.mem_bank[1336],db_even.mem_bank[1336],db_odd.mem_bank[1337],db_even.mem_bank[1337],db_odd.mem_bank[1338],db_even.mem_bank[1338],db_odd.mem_bank[1339],db_even.mem_bank[1339],db_odd.mem_bank[1340],db_even.mem_bank[1340],db_odd.mem_bank[1341],db_even.mem_bank[1341],db_odd.mem_bank[1342],db_even.mem_bank[1342],db_odd.mem_bank[1343],db_even.mem_bank[1343],db_odd.mem_bank[1344],db_even.mem_bank[1344],db_odd.mem_bank[1345],db_even.mem_bank[1345],db_odd.mem_bank[1346],db_even.mem_bank[1346],db_odd.mem_bank[1347],db_even.mem_bank[1347],db_odd.mem_bank[1348],db_even.mem_bank[1348],db_odd.mem_bank[1349],db_even.mem_bank[1349],db_odd.mem_bank[1350],db_even.mem_bank[1350],db_odd.mem_bank[1351],db_even.mem_bank[1351],db_odd.mem_bank[1352],db_even.mem_bank[1352],db_odd.mem_bank[1353],db_even.mem_bank[1353],db_odd.mem_bank[1354],db_even.mem_bank[1354],db_odd.mem_bank[1355],db_even.mem_bank[1355],db_odd.mem_bank[1356],db_even.mem_bank[1356],db_odd.mem_bank[1357],db_even.mem_bank[1357],db_odd.mem_bank[1358],db_even.mem_bank[1358],db_odd.mem_bank[1359],db_even.mem_bank[1359],db_odd.mem_bank[1360],db_even.mem_bank[1360],db_odd.mem_bank[1361],db_even.mem_bank[1361],db_odd.mem_bank[1362],db_even.mem_bank[1362],db_odd.mem_bank[1363],db_even.mem_bank[1363],db_odd.mem_bank[1364],db_even.mem_bank[1364],db_odd.mem_bank[1365],db_even.mem_bank[1365],db_odd.mem_bank[1366],db_even.mem_bank[1366],db_odd.mem_bank[1367],db_even.mem_bank[1367],db_odd.mem_bank[1368],db_even.mem_bank[1368],db_odd.mem_bank[1369],db_even.mem_bank[1369],db_odd.mem_bank[1370],db_even.mem_bank[1370],db_odd.mem_bank[1371],db_even.mem_bank[1371],db_odd.mem_bank[1372],db_even.mem_bank[1372],db_odd.mem_bank[1373],db_even.mem_bank[1373],db_odd.mem_bank[1374],db_even.mem_bank[1374],db_odd.mem_bank[1375],db_even.mem_bank[1375],db_odd.mem_bank[1376],db_even.mem_bank[1376],db_odd.mem_bank[1377],db_even.mem_bank[1377],db_odd.mem_bank[1378],db_even.mem_bank[1378],db_odd.mem_bank[1379],db_even.mem_bank[1379],db_odd.mem_bank[1380],db_even.mem_bank[1380],db_odd.mem_bank[1381],db_even.mem_bank[1381],db_odd.mem_bank[1382],db_even.mem_bank[1382],db_odd.mem_bank[1383],db_even.mem_bank[1383],db_odd.mem_bank[1384],db_even.mem_bank[1384],db_odd.mem_bank[1385],db_even.mem_bank[1385],db_odd.mem_bank[1386],db_even.mem_bank[1386],db_odd.mem_bank[1387],db_even.mem_bank[1387],db_odd.mem_bank[1388],db_even.mem_bank[1388],db_odd.mem_bank[1389],db_even.mem_bank[1389],db_odd.mem_bank[1390],db_even.mem_bank[1390],db_odd.mem_bank[1391],db_even.mem_bank[1391],db_odd.mem_bank[1392],db_even.mem_bank[1392],db_odd.mem_bank[1393],db_even.mem_bank[1393],db_odd.mem_bank[1394],db_even.mem_bank[1394],db_odd.mem_bank[1395],db_even.mem_bank[1395],db_odd.mem_bank[1396],db_even.mem_bank[1396],db_odd.mem_bank[1397],db_even.mem_bank[1397],db_odd.mem_bank[1398],db_even.mem_bank[1398],db_odd.mem_bank[1399],db_even.mem_bank[1399],db_odd.mem_bank[1400],db_even.mem_bank[1400],db_odd.mem_bank[1401],db_even.mem_bank[1401],db_odd.mem_bank[1402],db_even.mem_bank[1402],db_odd.mem_bank[1403],db_even.mem_bank[1403],db_odd.mem_bank[1404],db_even.mem_bank[1404],db_odd.mem_bank[1405],db_even.mem_bank[1405],db_odd.mem_bank[1406],db_even.mem_bank[1406],db_odd.mem_bank[1407],db_even.mem_bank[1407],db_odd.mem_bank[1408],db_even.mem_bank[1408],db_odd.mem_bank[1409],db_even.mem_bank[1409],db_odd.mem_bank[1410],db_even.mem_bank[1410],db_odd.mem_bank[1411],db_even.mem_bank[1411],db_odd.mem_bank[1412],db_even.mem_bank[1412],db_odd.mem_bank[1413],db_even.mem_bank[1413],db_odd.mem_bank[1414],db_even.mem_bank[1414],db_odd.mem_bank[1415],db_even.mem_bank[1415],db_odd.mem_bank[1416],db_even.mem_bank[1416],db_odd.mem_bank[1417],db_even.mem_bank[1417],db_odd.mem_bank[1418],db_even.mem_bank[1418],db_odd.mem_bank[1419],db_even.mem_bank[1419],db_odd.mem_bank[1420],db_even.mem_bank[1420],db_odd.mem_bank[1421],db_even.mem_bank[1421],db_odd.mem_bank[1422],db_even.mem_bank[1422],db_odd.mem_bank[1423],db_even.mem_bank[1423],db_odd.mem_bank[1424],db_even.mem_bank[1424],db_odd.mem_bank[1425],db_even.mem_bank[1425],db_odd.mem_bank[1426],db_even.mem_bank[1426],db_odd.mem_bank[1427],db_even.mem_bank[1427],db_odd.mem_bank[1428],db_even.mem_bank[1428],db_odd.mem_bank[1429],db_even.mem_bank[1429],db_odd.mem_bank[1430],db_even.mem_bank[1430],db_odd.mem_bank[1431],db_even.mem_bank[1431],db_odd.mem_bank[1432],db_even.mem_bank[1432],db_odd.mem_bank[1433],db_even.mem_bank[1433],db_odd.mem_bank[1434],db_even.mem_bank[1434],db_odd.mem_bank[1435],db_even.mem_bank[1435],db_odd.mem_bank[1436],db_even.mem_bank[1436],db_odd.mem_bank[1437],db_even.mem_bank[1437],db_odd.mem_bank[1438],db_even.mem_bank[1438],db_odd.mem_bank[1439],db_even.mem_bank[1439],db_odd.mem_bank[1440],db_even.mem_bank[1440],db_odd.mem_bank[1441],db_even.mem_bank[1441],db_odd.mem_bank[1442],db_even.mem_bank[1442],db_odd.mem_bank[1443],db_even.mem_bank[1443],db_odd.mem_bank[1444],db_even.mem_bank[1444],db_odd.mem_bank[1445],db_even.mem_bank[1445],db_odd.mem_bank[1446],db_even.mem_bank[1446],db_odd.mem_bank[1447],db_even.mem_bank[1447],db_odd.mem_bank[1448],db_even.mem_bank[1448],db_odd.mem_bank[1449],db_even.mem_bank[1449],db_odd.mem_bank[1450],db_even.mem_bank[1450],db_odd.mem_bank[1451],db_even.mem_bank[1451],db_odd.mem_bank[1452],db_even.mem_bank[1452],db_odd.mem_bank[1453],db_even.mem_bank[1453],db_odd.mem_bank[1454],db_even.mem_bank[1454],db_odd.mem_bank[1455],db_even.mem_bank[1455],db_odd.mem_bank[1456],db_even.mem_bank[1456],db_odd.mem_bank[1457],db_even.mem_bank[1457],db_odd.mem_bank[1458],db_even.mem_bank[1458],db_odd.mem_bank[1459],db_even.mem_bank[1459],db_odd.mem_bank[1460],db_even.mem_bank[1460],db_odd.mem_bank[1461],db_even.mem_bank[1461],db_odd.mem_bank[1462],db_even.mem_bank[1462],db_odd.mem_bank[1463],db_even.mem_bank[1463],db_odd.mem_bank[1464],db_even.mem_bank[1464],db_odd.mem_bank[1465],db_even.mem_bank[1465],db_odd.mem_bank[1466],db_even.mem_bank[1466],db_odd.mem_bank[1467],db_even.mem_bank[1467],db_odd.mem_bank[1468],db_even.mem_bank[1468],db_odd.mem_bank[1469],db_even.mem_bank[1469],db_odd.mem_bank[1470],db_even.mem_bank[1470],db_odd.mem_bank[1471],db_even.mem_bank[1471],db_odd.mem_bank[1472],db_even.mem_bank[1472],db_odd.mem_bank[1473],db_even.mem_bank[1473],db_odd.mem_bank[1474],db_even.mem_bank[1474],db_odd.mem_bank[1475],db_even.mem_bank[1475],db_odd.mem_bank[1476],db_even.mem_bank[1476],db_odd.mem_bank[1477],db_even.mem_bank[1477],db_odd.mem_bank[1478],db_even.mem_bank[1478],db_odd.mem_bank[1479],db_even.mem_bank[1479],db_odd.mem_bank[1480],db_even.mem_bank[1480],db_odd.mem_bank[1481],db_even.mem_bank[1481],db_odd.mem_bank[1482],db_even.mem_bank[1482],db_odd.mem_bank[1483],db_even.mem_bank[1483],db_odd.mem_bank[1484],db_even.mem_bank[1484],db_odd.mem_bank[1485],db_even.mem_bank[1485],db_odd.mem_bank[1486],db_even.mem_bank[1486],db_odd.mem_bank[1487],db_even.mem_bank[1487],db_odd.mem_bank[1488],db_even.mem_bank[1488],db_odd.mem_bank[1489],db_even.mem_bank[1489],db_odd.mem_bank[1490],db_even.mem_bank[1490],db_odd.mem_bank[1491],db_even.mem_bank[1491],db_odd.mem_bank[1492],db_even.mem_bank[1492],db_odd.mem_bank[1493],db_even.mem_bank[1493],db_odd.mem_bank[1494],db_even.mem_bank[1494],db_odd.mem_bank[1495],db_even.mem_bank[1495],db_odd.mem_bank[1496],db_even.mem_bank[1496],db_odd.mem_bank[1497],db_even.mem_bank[1497],db_odd.mem_bank[1498],db_even.mem_bank[1498],db_odd.mem_bank[1499],db_even.mem_bank[1499],db_odd.mem_bank[1500],db_even.mem_bank[1500],db_odd.mem_bank[1501],db_even.mem_bank[1501],db_odd.mem_bank[1502],db_even.mem_bank[1502],db_odd.mem_bank[1503],db_even.mem_bank[1503],db_odd.mem_bank[1504],db_even.mem_bank[1504],db_odd.mem_bank[1505],db_even.mem_bank[1505],db_odd.mem_bank[1506],db_even.mem_bank[1506],db_odd.mem_bank[1507],db_even.mem_bank[1507],db_odd.mem_bank[1508],db_even.mem_bank[1508],db_odd.mem_bank[1509],db_even.mem_bank[1509],db_odd.mem_bank[1510],db_even.mem_bank[1510],db_odd.mem_bank[1511],db_even.mem_bank[1511],db_odd.mem_bank[1512],db_even.mem_bank[1512],db_odd.mem_bank[1513],db_even.mem_bank[1513],db_odd.mem_bank[1514],db_even.mem_bank[1514],db_odd.mem_bank[1515],db_even.mem_bank[1515],db_odd.mem_bank[1516],db_even.mem_bank[1516],db_odd.mem_bank[1517],db_even.mem_bank[1517],db_odd.mem_bank[1518],db_even.mem_bank[1518],db_odd.mem_bank[1519],db_even.mem_bank[1519],db_odd.mem_bank[1520],db_even.mem_bank[1520],db_odd.mem_bank[1521],db_even.mem_bank[1521],db_odd.mem_bank[1522],db_even.mem_bank[1522],db_odd.mem_bank[1523],db_even.mem_bank[1523],db_odd.mem_bank[1524],db_even.mem_bank[1524],db_odd.mem_bank[1525],db_even.mem_bank[1525],db_odd.mem_bank[1526],db_even.mem_bank[1526],db_odd.mem_bank[1527],db_even.mem_bank[1527],db_odd.mem_bank[1528],db_even.mem_bank[1528],db_odd.mem_bank[1529],db_even.mem_bank[1529],db_odd.mem_bank[1530],db_even.mem_bank[1530],db_odd.mem_bank[1531],db_even.mem_bank[1531],db_odd.mem_bank[1532],db_even.mem_bank[1532],db_odd.mem_bank[1533],db_even.mem_bank[1533],db_odd.mem_bank[1534],db_even.mem_bank[1534],db_odd.mem_bank[1535],db_even.mem_bank[1535],db_odd.mem_bank[1536],db_even.mem_bank[1536],db_odd.mem_bank[1537],db_even.mem_bank[1537],db_odd.mem_bank[1538],db_even.mem_bank[1538],db_odd.mem_bank[1539],db_even.mem_bank[1539],db_odd.mem_bank[1540],db_even.mem_bank[1540],db_odd.mem_bank[1541],db_even.mem_bank[1541],db_odd.mem_bank[1542],db_even.mem_bank[1542],db_odd.mem_bank[1543],db_even.mem_bank[1543],db_odd.mem_bank[1544],db_even.mem_bank[1544],db_odd.mem_bank[1545],db_even.mem_bank[1545],db_odd.mem_bank[1546],db_even.mem_bank[1546],db_odd.mem_bank[1547],db_even.mem_bank[1547],db_odd.mem_bank[1548],db_even.mem_bank[1548],db_odd.mem_bank[1549],db_even.mem_bank[1549],db_odd.mem_bank[1550],db_even.mem_bank[1550],db_odd.mem_bank[1551],db_even.mem_bank[1551],db_odd.mem_bank[1552],db_even.mem_bank[1552],db_odd.mem_bank[1553],db_even.mem_bank[1553],db_odd.mem_bank[1554],db_even.mem_bank[1554],db_odd.mem_bank[1555],db_even.mem_bank[1555],db_odd.mem_bank[1556],db_even.mem_bank[1556],db_odd.mem_bank[1557],db_even.mem_bank[1557],db_odd.mem_bank[1558],db_even.mem_bank[1558],db_odd.mem_bank[1559],db_even.mem_bank[1559],db_odd.mem_bank[1560],db_even.mem_bank[1560],db_odd.mem_bank[1561],db_even.mem_bank[1561],db_odd.mem_bank[1562],db_even.mem_bank[1562],db_odd.mem_bank[1563],db_even.mem_bank[1563],db_odd.mem_bank[1564],db_even.mem_bank[1564],db_odd.mem_bank[1565],db_even.mem_bank[1565],db_odd.mem_bank[1566],db_even.mem_bank[1566],db_odd.mem_bank[1567],db_even.mem_bank[1567],db_odd.mem_bank[1568],db_even.mem_bank[1568],db_odd.mem_bank[1569],db_even.mem_bank[1569],db_odd.mem_bank[1570],db_even.mem_bank[1570],db_odd.mem_bank[1571],db_even.mem_bank[1571],db_odd.mem_bank[1572],db_even.mem_bank[1572],db_odd.mem_bank[1573],db_even.mem_bank[1573],db_odd.mem_bank[1574],db_even.mem_bank[1574],db_odd.mem_bank[1575],db_even.mem_bank[1575],db_odd.mem_bank[1576],db_even.mem_bank[1576],db_odd.mem_bank[1577],db_even.mem_bank[1577],db_odd.mem_bank[1578],db_even.mem_bank[1578],db_odd.mem_bank[1579],db_even.mem_bank[1579],db_odd.mem_bank[1580],db_even.mem_bank[1580],db_odd.mem_bank[1581],db_even.mem_bank[1581],db_odd.mem_bank[1582],db_even.mem_bank[1582],db_odd.mem_bank[1583],db_even.mem_bank[1583],db_odd.mem_bank[1584],db_even.mem_bank[1584],db_odd.mem_bank[1585],db_even.mem_bank[1585],db_odd.mem_bank[1586],db_even.mem_bank[1586],db_odd.mem_bank[1587],db_even.mem_bank[1587],db_odd.mem_bank[1588],db_even.mem_bank[1588],db_odd.mem_bank[1589],db_even.mem_bank[1589],db_odd.mem_bank[1590],db_even.mem_bank[1590],db_odd.mem_bank[1591],db_even.mem_bank[1591],db_odd.mem_bank[1592],db_even.mem_bank[1592],db_odd.mem_bank[1593],db_even.mem_bank[1593],db_odd.mem_bank[1594],db_even.mem_bank[1594],db_odd.mem_bank[1595],db_even.mem_bank[1595],db_odd.mem_bank[1596],db_even.mem_bank[1596],db_odd.mem_bank[1597],db_even.mem_bank[1597],db_odd.mem_bank[1598],db_even.mem_bank[1598],db_odd.mem_bank[1599],db_even.mem_bank[1599],db_odd.mem_bank[1600],db_even.mem_bank[1600],db_odd.mem_bank[1601],db_even.mem_bank[1601],db_odd.mem_bank[1602],db_even.mem_bank[1602],db_odd.mem_bank[1603],db_even.mem_bank[1603],db_odd.mem_bank[1604],db_even.mem_bank[1604],db_odd.mem_bank[1605],db_even.mem_bank[1605],db_odd.mem_bank[1606],db_even.mem_bank[1606],db_odd.mem_bank[1607],db_even.mem_bank[1607],db_odd.mem_bank[1608],db_even.mem_bank[1608],db_odd.mem_bank[1609],db_even.mem_bank[1609],db_odd.mem_bank[1610],db_even.mem_bank[1610],db_odd.mem_bank[1611],db_even.mem_bank[1611],db_odd.mem_bank[1612],db_even.mem_bank[1612],db_odd.mem_bank[1613],db_even.mem_bank[1613],db_odd.mem_bank[1614],db_even.mem_bank[1614],db_odd.mem_bank[1615],db_even.mem_bank[1615],db_odd.mem_bank[1616],db_even.mem_bank[1616],db_odd.mem_bank[1617],db_even.mem_bank[1617],db_odd.mem_bank[1618],db_even.mem_bank[1618],db_odd.mem_bank[1619],db_even.mem_bank[1619],db_odd.mem_bank[1620],db_even.mem_bank[1620],db_odd.mem_bank[1621],db_even.mem_bank[1621],db_odd.mem_bank[1622],db_even.mem_bank[1622],db_odd.mem_bank[1623],db_even.mem_bank[1623],db_odd.mem_bank[1624],db_even.mem_bank[1624],db_odd.mem_bank[1625],db_even.mem_bank[1625],db_odd.mem_bank[1626],db_even.mem_bank[1626],db_odd.mem_bank[1627],db_even.mem_bank[1627],db_odd.mem_bank[1628],db_even.mem_bank[1628],db_odd.mem_bank[1629],db_even.mem_bank[1629],db_odd.mem_bank[1630],db_even.mem_bank[1630],db_odd.mem_bank[1631],db_even.mem_bank[1631],db_odd.mem_bank[1632],db_even.mem_bank[1632],db_odd.mem_bank[1633],db_even.mem_bank[1633],db_odd.mem_bank[1634],db_even.mem_bank[1634],db_odd.mem_bank[1635],db_even.mem_bank[1635],db_odd.mem_bank[1636],db_even.mem_bank[1636],db_odd.mem_bank[1637],db_even.mem_bank[1637],db_odd.mem_bank[1638],db_even.mem_bank[1638],db_odd.mem_bank[1639],db_even.mem_bank[1639],db_odd.mem_bank[1640],db_even.mem_bank[1640],db_odd.mem_bank[1641],db_even.mem_bank[1641],db_odd.mem_bank[1642],db_even.mem_bank[1642],db_odd.mem_bank[1643],db_even.mem_bank[1643],db_odd.mem_bank[1644],db_even.mem_bank[1644],db_odd.mem_bank[1645],db_even.mem_bank[1645],db_odd.mem_bank[1646],db_even.mem_bank[1646],db_odd.mem_bank[1647],db_even.mem_bank[1647],db_odd.mem_bank[1648],db_even.mem_bank[1648],db_odd.mem_bank[1649],db_even.mem_bank[1649],db_odd.mem_bank[1650],db_even.mem_bank[1650],db_odd.mem_bank[1651],db_even.mem_bank[1651],db_odd.mem_bank[1652],db_even.mem_bank[1652],db_odd.mem_bank[1653],db_even.mem_bank[1653],db_odd.mem_bank[1654],db_even.mem_bank[1654],db_odd.mem_bank[1655],db_even.mem_bank[1655],db_odd.mem_bank[1656],db_even.mem_bank[1656],db_odd.mem_bank[1657],db_even.mem_bank[1657],db_odd.mem_bank[1658],db_even.mem_bank[1658],db_odd.mem_bank[1659],db_even.mem_bank[1659],db_odd.mem_bank[1660],db_even.mem_bank[1660],db_odd.mem_bank[1661],db_even.mem_bank[1661],db_odd.mem_bank[1662],db_even.mem_bank[1662],db_odd.mem_bank[1663],db_even.mem_bank[1663],db_odd.mem_bank[1664],db_even.mem_bank[1664],db_odd.mem_bank[1665],db_even.mem_bank[1665],db_odd.mem_bank[1666],db_even.mem_bank[1666],db_odd.mem_bank[1667],db_even.mem_bank[1667],db_odd.mem_bank[1668],db_even.mem_bank[1668],db_odd.mem_bank[1669],db_even.mem_bank[1669],db_odd.mem_bank[1670],db_even.mem_bank[1670],db_odd.mem_bank[1671],db_even.mem_bank[1671],db_odd.mem_bank[1672],db_even.mem_bank[1672],db_odd.mem_bank[1673],db_even.mem_bank[1673],db_odd.mem_bank[1674],db_even.mem_bank[1674],db_odd.mem_bank[1675],db_even.mem_bank[1675],db_odd.mem_bank[1676],db_even.mem_bank[1676],db_odd.mem_bank[1677],db_even.mem_bank[1677],db_odd.mem_bank[1678],db_even.mem_bank[1678],db_odd.mem_bank[1679],db_even.mem_bank[1679],db_odd.mem_bank[1680],db_even.mem_bank[1680],db_odd.mem_bank[1681],db_even.mem_bank[1681],db_odd.mem_bank[1682],db_even.mem_bank[1682],db_odd.mem_bank[1683],db_even.mem_bank[1683],db_odd.mem_bank[1684],db_even.mem_bank[1684],db_odd.mem_bank[1685],db_even.mem_bank[1685],db_odd.mem_bank[1686],db_even.mem_bank[1686],db_odd.mem_bank[1687],db_even.mem_bank[1687],db_odd.mem_bank[1688],db_even.mem_bank[1688],db_odd.mem_bank[1689],db_even.mem_bank[1689],db_odd.mem_bank[1690],db_even.mem_bank[1690],db_odd.mem_bank[1691],db_even.mem_bank[1691],db_odd.mem_bank[1692],db_even.mem_bank[1692],db_odd.mem_bank[1693],db_even.mem_bank[1693],db_odd.mem_bank[1694],db_even.mem_bank[1694],db_odd.mem_bank[1695],db_even.mem_bank[1695],db_odd.mem_bank[1696],db_even.mem_bank[1696],db_odd.mem_bank[1697],db_even.mem_bank[1697],db_odd.mem_bank[1698],db_even.mem_bank[1698],db_odd.mem_bank[1699],db_even.mem_bank[1699],db_odd.mem_bank[1700],db_even.mem_bank[1700],db_odd.mem_bank[1701],db_even.mem_bank[1701],db_odd.mem_bank[1702],db_even.mem_bank[1702],db_odd.mem_bank[1703],db_even.mem_bank[1703],db_odd.mem_bank[1704],db_even.mem_bank[1704],db_odd.mem_bank[1705],db_even.mem_bank[1705],db_odd.mem_bank[1706],db_even.mem_bank[1706],db_odd.mem_bank[1707],db_even.mem_bank[1707],db_odd.mem_bank[1708],db_even.mem_bank[1708],db_odd.mem_bank[1709],db_even.mem_bank[1709],db_odd.mem_bank[1710],db_even.mem_bank[1710],db_odd.mem_bank[1711],db_even.mem_bank[1711],db_odd.mem_bank[1712],db_even.mem_bank[1712],db_odd.mem_bank[1713],db_even.mem_bank[1713],db_odd.mem_bank[1714],db_even.mem_bank[1714],db_odd.mem_bank[1715],db_even.mem_bank[1715],db_odd.mem_bank[1716],db_even.mem_bank[1716],db_odd.mem_bank[1717],db_even.mem_bank[1717],db_odd.mem_bank[1718],db_even.mem_bank[1718],db_odd.mem_bank[1719],db_even.mem_bank[1719],db_odd.mem_bank[1720],db_even.mem_bank[1720],db_odd.mem_bank[1721],db_even.mem_bank[1721],db_odd.mem_bank[1722],db_even.mem_bank[1722],db_odd.mem_bank[1723],db_even.mem_bank[1723],db_odd.mem_bank[1724],db_even.mem_bank[1724],db_odd.mem_bank[1725],db_even.mem_bank[1725],db_odd.mem_bank[1726],db_even.mem_bank[1726],db_odd.mem_bank[1727],db_even.mem_bank[1727],db_odd.mem_bank[1728],db_even.mem_bank[1728],db_odd.mem_bank[1729],db_even.mem_bank[1729],db_odd.mem_bank[1730],db_even.mem_bank[1730],db_odd.mem_bank[1731],db_even.mem_bank[1731],db_odd.mem_bank[1732],db_even.mem_bank[1732],db_odd.mem_bank[1733],db_even.mem_bank[1733],db_odd.mem_bank[1734],db_even.mem_bank[1734],db_odd.mem_bank[1735],db_even.mem_bank[1735],db_odd.mem_bank[1736],db_even.mem_bank[1736],db_odd.mem_bank[1737],db_even.mem_bank[1737],db_odd.mem_bank[1738],db_even.mem_bank[1738],db_odd.mem_bank[1739],db_even.mem_bank[1739],db_odd.mem_bank[1740],db_even.mem_bank[1740],db_odd.mem_bank[1741],db_even.mem_bank[1741],db_odd.mem_bank[1742],db_even.mem_bank[1742],db_odd.mem_bank[1743],db_even.mem_bank[1743],db_odd.mem_bank[1744],db_even.mem_bank[1744],db_odd.mem_bank[1745],db_even.mem_bank[1745],db_odd.mem_bank[1746],db_even.mem_bank[1746],db_odd.mem_bank[1747],db_even.mem_bank[1747],db_odd.mem_bank[1748],db_even.mem_bank[1748],db_odd.mem_bank[1749],db_even.mem_bank[1749],db_odd.mem_bank[1750],db_even.mem_bank[1750],db_odd.mem_bank[1751],db_even.mem_bank[1751],db_odd.mem_bank[1752],db_even.mem_bank[1752],db_odd.mem_bank[1753],db_even.mem_bank[1753],db_odd.mem_bank[1754],db_even.mem_bank[1754],db_odd.mem_bank[1755],db_even.mem_bank[1755],db_odd.mem_bank[1756],db_even.mem_bank[1756],db_odd.mem_bank[1757],db_even.mem_bank[1757],db_odd.mem_bank[1758],db_even.mem_bank[1758],db_odd.mem_bank[1759],db_even.mem_bank[1759],db_odd.mem_bank[1760],db_even.mem_bank[1760],db_odd.mem_bank[1761],db_even.mem_bank[1761],db_odd.mem_bank[1762],db_even.mem_bank[1762],db_odd.mem_bank[1763],db_even.mem_bank[1763],db_odd.mem_bank[1764],db_even.mem_bank[1764],db_odd.mem_bank[1765],db_even.mem_bank[1765],db_odd.mem_bank[1766],db_even.mem_bank[1766],db_odd.mem_bank[1767],db_even.mem_bank[1767],db_odd.mem_bank[1768],db_even.mem_bank[1768],db_odd.mem_bank[1769],db_even.mem_bank[1769],db_odd.mem_bank[1770],db_even.mem_bank[1770],db_odd.mem_bank[1771],db_even.mem_bank[1771],db_odd.mem_bank[1772],db_even.mem_bank[1772],db_odd.mem_bank[1773],db_even.mem_bank[1773],db_odd.mem_bank[1774],db_even.mem_bank[1774],db_odd.mem_bank[1775],db_even.mem_bank[1775],db_odd.mem_bank[1776],db_even.mem_bank[1776],db_odd.mem_bank[1777],db_even.mem_bank[1777],db_odd.mem_bank[1778],db_even.mem_bank[1778],db_odd.mem_bank[1779],db_even.mem_bank[1779],db_odd.mem_bank[1780],db_even.mem_bank[1780],db_odd.mem_bank[1781],db_even.mem_bank[1781],db_odd.mem_bank[1782],db_even.mem_bank[1782],db_odd.mem_bank[1783],db_even.mem_bank[1783],db_odd.mem_bank[1784],db_even.mem_bank[1784],db_odd.mem_bank[1785],db_even.mem_bank[1785],db_odd.mem_bank[1786],db_even.mem_bank[1786],db_odd.mem_bank[1787],db_even.mem_bank[1787],db_odd.mem_bank[1788],db_even.mem_bank[1788],db_odd.mem_bank[1789],db_even.mem_bank[1789],db_odd.mem_bank[1790],db_even.mem_bank[1790],db_odd.mem_bank[1791],db_even.mem_bank[1791],db_odd.mem_bank[1792],db_even.mem_bank[1792],db_odd.mem_bank[1793],db_even.mem_bank[1793],db_odd.mem_bank[1794],db_even.mem_bank[1794],db_odd.mem_bank[1795],db_even.mem_bank[1795],db_odd.mem_bank[1796],db_even.mem_bank[1796],db_odd.mem_bank[1797],db_even.mem_bank[1797],db_odd.mem_bank[1798],db_even.mem_bank[1798],db_odd.mem_bank[1799],db_even.mem_bank[1799],db_odd.mem_bank[1800],db_even.mem_bank[1800],db_odd.mem_bank[1801],db_even.mem_bank[1801],db_odd.mem_bank[1802],db_even.mem_bank[1802],db_odd.mem_bank[1803],db_even.mem_bank[1803],db_odd.mem_bank[1804],db_even.mem_bank[1804],db_odd.mem_bank[1805],db_even.mem_bank[1805],db_odd.mem_bank[1806],db_even.mem_bank[1806],db_odd.mem_bank[1807],db_even.mem_bank[1807],db_odd.mem_bank[1808],db_even.mem_bank[1808],db_odd.mem_bank[1809],db_even.mem_bank[1809],db_odd.mem_bank[1810],db_even.mem_bank[1810],db_odd.mem_bank[1811],db_even.mem_bank[1811],db_odd.mem_bank[1812],db_even.mem_bank[1812],db_odd.mem_bank[1813],db_even.mem_bank[1813],db_odd.mem_bank[1814],db_even.mem_bank[1814],db_odd.mem_bank[1815],db_even.mem_bank[1815],db_odd.mem_bank[1816],db_even.mem_bank[1816],db_odd.mem_bank[1817],db_even.mem_bank[1817],db_odd.mem_bank[1818],db_even.mem_bank[1818],db_odd.mem_bank[1819],db_even.mem_bank[1819],db_odd.mem_bank[1820],db_even.mem_bank[1820],db_odd.mem_bank[1821],db_even.mem_bank[1821],db_odd.mem_bank[1822],db_even.mem_bank[1822],db_odd.mem_bank[1823],db_even.mem_bank[1823],db_odd.mem_bank[1824],db_even.mem_bank[1824],db_odd.mem_bank[1825],db_even.mem_bank[1825],db_odd.mem_bank[1826],db_even.mem_bank[1826],db_odd.mem_bank[1827],db_even.mem_bank[1827],db_odd.mem_bank[1828],db_even.mem_bank[1828],db_odd.mem_bank[1829],db_even.mem_bank[1829],db_odd.mem_bank[1830],db_even.mem_bank[1830],db_odd.mem_bank[1831],db_even.mem_bank[1831],db_odd.mem_bank[1832],db_even.mem_bank[1832],db_odd.mem_bank[1833],db_even.mem_bank[1833],db_odd.mem_bank[1834],db_even.mem_bank[1834],db_odd.mem_bank[1835],db_even.mem_bank[1835],db_odd.mem_bank[1836],db_even.mem_bank[1836],db_odd.mem_bank[1837],db_even.mem_bank[1837],db_odd.mem_bank[1838],db_even.mem_bank[1838],db_odd.mem_bank[1839],db_even.mem_bank[1839],db_odd.mem_bank[1840],db_even.mem_bank[1840],db_odd.mem_bank[1841],db_even.mem_bank[1841],db_odd.mem_bank[1842],db_even.mem_bank[1842],db_odd.mem_bank[1843],db_even.mem_bank[1843],db_odd.mem_bank[1844],db_even.mem_bank[1844],db_odd.mem_bank[1845],db_even.mem_bank[1845],db_odd.mem_bank[1846],db_even.mem_bank[1846],db_odd.mem_bank[1847],db_even.mem_bank[1847],db_odd.mem_bank[1848],db_even.mem_bank[1848],db_odd.mem_bank[1849],db_even.mem_bank[1849],db_odd.mem_bank[1850],db_even.mem_bank[1850],db_odd.mem_bank[1851],db_even.mem_bank[1851],db_odd.mem_bank[1852],db_even.mem_bank[1852],db_odd.mem_bank[1853],db_even.mem_bank[1853],db_odd.mem_bank[1854],db_even.mem_bank[1854],db_odd.mem_bank[1855],db_even.mem_bank[1855],db_odd.mem_bank[1856],db_even.mem_bank[1856],db_odd.mem_bank[1857],db_even.mem_bank[1857],db_odd.mem_bank[1858],db_even.mem_bank[1858],db_odd.mem_bank[1859],db_even.mem_bank[1859],db_odd.mem_bank[1860],db_even.mem_bank[1860],db_odd.mem_bank[1861],db_even.mem_bank[1861],db_odd.mem_bank[1862],db_even.mem_bank[1862],db_odd.mem_bank[1863],db_even.mem_bank[1863],db_odd.mem_bank[1864],db_even.mem_bank[1864],db_odd.mem_bank[1865],db_even.mem_bank[1865],db_odd.mem_bank[1866],db_even.mem_bank[1866],db_odd.mem_bank[1867],db_even.mem_bank[1867],db_odd.mem_bank[1868],db_even.mem_bank[1868],db_odd.mem_bank[1869],db_even.mem_bank[1869],db_odd.mem_bank[1870],db_even.mem_bank[1870],db_odd.mem_bank[1871],db_even.mem_bank[1871],db_odd.mem_bank[1872],db_even.mem_bank[1872],db_odd.mem_bank[1873],db_even.mem_bank[1873],db_odd.mem_bank[1874],db_even.mem_bank[1874],db_odd.mem_bank[1875],db_even.mem_bank[1875],db_odd.mem_bank[1876],db_even.mem_bank[1876],db_odd.mem_bank[1877],db_even.mem_bank[1877],db_odd.mem_bank[1878],db_even.mem_bank[1878],db_odd.mem_bank[1879],db_even.mem_bank[1879],db_odd.mem_bank[1880],db_even.mem_bank[1880],db_odd.mem_bank[1881],db_even.mem_bank[1881],db_odd.mem_bank[1882],db_even.mem_bank[1882],db_odd.mem_bank[1883],db_even.mem_bank[1883],db_odd.mem_bank[1884],db_even.mem_bank[1884],db_odd.mem_bank[1885],db_even.mem_bank[1885],db_odd.mem_bank[1886],db_even.mem_bank[1886],db_odd.mem_bank[1887],db_even.mem_bank[1887],db_odd.mem_bank[1888],db_even.mem_bank[1888],db_odd.mem_bank[1889],db_even.mem_bank[1889],db_odd.mem_bank[1890],db_even.mem_bank[1890],db_odd.mem_bank[1891],db_even.mem_bank[1891],db_odd.mem_bank[1892],db_even.mem_bank[1892],db_odd.mem_bank[1893],db_even.mem_bank[1893],db_odd.mem_bank[1894],db_even.mem_bank[1894],db_odd.mem_bank[1895],db_even.mem_bank[1895],db_odd.mem_bank[1896],db_even.mem_bank[1896],db_odd.mem_bank[1897],db_even.mem_bank[1897],db_odd.mem_bank[1898],db_even.mem_bank[1898],db_odd.mem_bank[1899],db_even.mem_bank[1899],db_odd.mem_bank[1900],db_even.mem_bank[1900],db_odd.mem_bank[1901],db_even.mem_bank[1901],db_odd.mem_bank[1902],db_even.mem_bank[1902],db_odd.mem_bank[1903],db_even.mem_bank[1903],db_odd.mem_bank[1904],db_even.mem_bank[1904],db_odd.mem_bank[1905],db_even.mem_bank[1905],db_odd.mem_bank[1906],db_even.mem_bank[1906],db_odd.mem_bank[1907],db_even.mem_bank[1907],db_odd.mem_bank[1908],db_even.mem_bank[1908],db_odd.mem_bank[1909],db_even.mem_bank[1909],db_odd.mem_bank[1910],db_even.mem_bank[1910],db_odd.mem_bank[1911],db_even.mem_bank[1911],db_odd.mem_bank[1912],db_even.mem_bank[1912],db_odd.mem_bank[1913],db_even.mem_bank[1913],db_odd.mem_bank[1914],db_even.mem_bank[1914],db_odd.mem_bank[1915],db_even.mem_bank[1915],db_odd.mem_bank[1916],db_even.mem_bank[1916],db_odd.mem_bank[1917],db_even.mem_bank[1917],db_odd.mem_bank[1918],db_even.mem_bank[1918],db_odd.mem_bank[1919],db_even.mem_bank[1919],db_odd.mem_bank[1920],db_even.mem_bank[1920],db_odd.mem_bank[1921],db_even.mem_bank[1921],db_odd.mem_bank[1922],db_even.mem_bank[1922],db_odd.mem_bank[1923],db_even.mem_bank[1923],db_odd.mem_bank[1924],db_even.mem_bank[1924],db_odd.mem_bank[1925],db_even.mem_bank[1925],db_odd.mem_bank[1926],db_even.mem_bank[1926],db_odd.mem_bank[1927],db_even.mem_bank[1927],db_odd.mem_bank[1928],db_even.mem_bank[1928],db_odd.mem_bank[1929],db_even.mem_bank[1929],db_odd.mem_bank[1930],db_even.mem_bank[1930],db_odd.mem_bank[1931],db_even.mem_bank[1931],db_odd.mem_bank[1932],db_even.mem_bank[1932],db_odd.mem_bank[1933],db_even.mem_bank[1933],db_odd.mem_bank[1934],db_even.mem_bank[1934],db_odd.mem_bank[1935],db_even.mem_bank[1935],db_odd.mem_bank[1936],db_even.mem_bank[1936],db_odd.mem_bank[1937],db_even.mem_bank[1937],db_odd.mem_bank[1938],db_even.mem_bank[1938],db_odd.mem_bank[1939],db_even.mem_bank[1939],db_odd.mem_bank[1940],db_even.mem_bank[1940],db_odd.mem_bank[1941],db_even.mem_bank[1941],db_odd.mem_bank[1942],db_even.mem_bank[1942],db_odd.mem_bank[1943],db_even.mem_bank[1943],db_odd.mem_bank[1944],db_even.mem_bank[1944],db_odd.mem_bank[1945],db_even.mem_bank[1945],db_odd.mem_bank[1946],db_even.mem_bank[1946],db_odd.mem_bank[1947],db_even.mem_bank[1947],db_odd.mem_bank[1948],db_even.mem_bank[1948],db_odd.mem_bank[1949],db_even.mem_bank[1949],db_odd.mem_bank[1950],db_even.mem_bank[1950],db_odd.mem_bank[1951],db_even.mem_bank[1951],db_odd.mem_bank[1952],db_even.mem_bank[1952],db_odd.mem_bank[1953],db_even.mem_bank[1953],db_odd.mem_bank[1954],db_even.mem_bank[1954],db_odd.mem_bank[1955],db_even.mem_bank[1955],db_odd.mem_bank[1956],db_even.mem_bank[1956],db_odd.mem_bank[1957],db_even.mem_bank[1957],db_odd.mem_bank[1958],db_even.mem_bank[1958],db_odd.mem_bank[1959],db_even.mem_bank[1959],db_odd.mem_bank[1960],db_even.mem_bank[1960],db_odd.mem_bank[1961],db_even.mem_bank[1961],db_odd.mem_bank[1962],db_even.mem_bank[1962],db_odd.mem_bank[1963],db_even.mem_bank[1963],db_odd.mem_bank[1964],db_even.mem_bank[1964],db_odd.mem_bank[1965],db_even.mem_bank[1965],db_odd.mem_bank[1966],db_even.mem_bank[1966],db_odd.mem_bank[1967],db_even.mem_bank[1967],db_odd.mem_bank[1968],db_even.mem_bank[1968],db_odd.mem_bank[1969],db_even.mem_bank[1969],db_odd.mem_bank[1970],db_even.mem_bank[1970],db_odd.mem_bank[1971],db_even.mem_bank[1971],db_odd.mem_bank[1972],db_even.mem_bank[1972],db_odd.mem_bank[1973],db_even.mem_bank[1973],db_odd.mem_bank[1974],db_even.mem_bank[1974],db_odd.mem_bank[1975],db_even.mem_bank[1975],db_odd.mem_bank[1976],db_even.mem_bank[1976],db_odd.mem_bank[1977],db_even.mem_bank[1977],db_odd.mem_bank[1978],db_even.mem_bank[1978],db_odd.mem_bank[1979],db_even.mem_bank[1979],db_odd.mem_bank[1980],db_even.mem_bank[1980],db_odd.mem_bank[1981],db_even.mem_bank[1981],db_odd.mem_bank[1982],db_even.mem_bank[1982],db_odd.mem_bank[1983],db_even.mem_bank[1983],db_odd.mem_bank[1984],db_even.mem_bank[1984],db_odd.mem_bank[1985],db_even.mem_bank[1985],db_odd.mem_bank[1986],db_even.mem_bank[1986],db_odd.mem_bank[1987],db_even.mem_bank[1987],db_odd.mem_bank[1988],db_even.mem_bank[1988],db_odd.mem_bank[1989],db_even.mem_bank[1989],db_odd.mem_bank[1990],db_even.mem_bank[1990],db_odd.mem_bank[1991],db_even.mem_bank[1991],db_odd.mem_bank[1992],db_even.mem_bank[1992],db_odd.mem_bank[1993],db_even.mem_bank[1993],db_odd.mem_bank[1994],db_even.mem_bank[1994],db_odd.mem_bank[1995],db_even.mem_bank[1995],db_odd.mem_bank[1996],db_even.mem_bank[1996],db_odd.mem_bank[1997],db_even.mem_bank[1997],db_odd.mem_bank[1998],db_even.mem_bank[1998],db_odd.mem_bank[1999],db_even.mem_bank[1999],db_odd.mem_bank[2000],db_even.mem_bank[2000],db_odd.mem_bank[2001],db_even.mem_bank[2001],db_odd.mem_bank[2002],db_even.mem_bank[2002],db_odd.mem_bank[2003],db_even.mem_bank[2003],db_odd.mem_bank[2004],db_even.mem_bank[2004],db_odd.mem_bank[2005],db_even.mem_bank[2005],db_odd.mem_bank[2006],db_even.mem_bank[2006],db_odd.mem_bank[2007],db_even.mem_bank[2007],db_odd.mem_bank[2008],db_even.mem_bank[2008],db_odd.mem_bank[2009],db_even.mem_bank[2009],db_odd.mem_bank[2010],db_even.mem_bank[2010],db_odd.mem_bank[2011],db_even.mem_bank[2011],db_odd.mem_bank[2012],db_even.mem_bank[2012],db_odd.mem_bank[2013],db_even.mem_bank[2013],db_odd.mem_bank[2014],db_even.mem_bank[2014],db_odd.mem_bank[2015],db_even.mem_bank[2015],db_odd.mem_bank[2016],db_even.mem_bank[2016],db_odd.mem_bank[2017],db_even.mem_bank[2017],db_odd.mem_bank[2018],db_even.mem_bank[2018],db_odd.mem_bank[2019],db_even.mem_bank[2019],db_odd.mem_bank[2020],db_even.mem_bank[2020],db_odd.mem_bank[2021],db_even.mem_bank[2021],db_odd.mem_bank[2022],db_even.mem_bank[2022],db_odd.mem_bank[2023],db_even.mem_bank[2023],db_odd.mem_bank[2024],db_even.mem_bank[2024],db_odd.mem_bank[2025],db_even.mem_bank[2025],db_odd.mem_bank[2026],db_even.mem_bank[2026],db_odd.mem_bank[2027],db_even.mem_bank[2027],db_odd.mem_bank[2028],db_even.mem_bank[2028],db_odd.mem_bank[2029],db_even.mem_bank[2029],db_odd.mem_bank[2030],db_even.mem_bank[2030],db_odd.mem_bank[2031],db_even.mem_bank[2031],db_odd.mem_bank[2032],db_even.mem_bank[2032],db_odd.mem_bank[2033],db_even.mem_bank[2033],db_odd.mem_bank[2034],db_even.mem_bank[2034],db_odd.mem_bank[2035],db_even.mem_bank[2035],db_odd.mem_bank[2036],db_even.mem_bank[2036],db_odd.mem_bank[2037],db_even.mem_bank[2037],db_odd.mem_bank[2038],db_even.mem_bank[2038],db_odd.mem_bank[2039],db_even.mem_bank[2039],db_odd.mem_bank[2040],db_even.mem_bank[2040],db_odd.mem_bank[2041],db_even.mem_bank[2041],db_odd.mem_bank[2042],db_even.mem_bank[2042],db_odd.mem_bank[2043],db_even.mem_bank[2043],db_odd.mem_bank[2044],db_even.mem_bank[2044],db_odd.mem_bank[2045],db_even.mem_bank[2045],db_odd.mem_bank[2046],db_even.mem_bank[2046],db_odd.mem_bank[2047],db_even.mem_bank[2047],db_odd.mem_bank[2048],db_even.mem_bank[2048],db_odd.mem_bank[2049],db_even.mem_bank[2049],db_odd.mem_bank[2050],db_even.mem_bank[2050],db_odd.mem_bank[2051],db_even.mem_bank[2051],db_odd.mem_bank[2052],db_even.mem_bank[2052],db_odd.mem_bank[2053],db_even.mem_bank[2053],db_odd.mem_bank[2054],db_even.mem_bank[2054],db_odd.mem_bank[2055],db_even.mem_bank[2055],db_odd.mem_bank[2056],db_even.mem_bank[2056],db_odd.mem_bank[2057],db_even.mem_bank[2057],db_odd.mem_bank[2058],db_even.mem_bank[2058],db_odd.mem_bank[2059],db_even.mem_bank[2059],db_odd.mem_bank[2060],db_even.mem_bank[2060],db_odd.mem_bank[2061],db_even.mem_bank[2061],db_odd.mem_bank[2062],db_even.mem_bank[2062],db_odd.mem_bank[2063],db_even.mem_bank[2063],db_odd.mem_bank[2064],db_even.mem_bank[2064],db_odd.mem_bank[2065],db_even.mem_bank[2065],db_odd.mem_bank[2066],db_even.mem_bank[2066],db_odd.mem_bank[2067],db_even.mem_bank[2067],db_odd.mem_bank[2068],db_even.mem_bank[2068],db_odd.mem_bank[2069],db_even.mem_bank[2069],db_odd.mem_bank[2070],db_even.mem_bank[2070],db_odd.mem_bank[2071],db_even.mem_bank[2071],db_odd.mem_bank[2072],db_even.mem_bank[2072],db_odd.mem_bank[2073],db_even.mem_bank[2073],db_odd.mem_bank[2074],db_even.mem_bank[2074],db_odd.mem_bank[2075],db_even.mem_bank[2075],db_odd.mem_bank[2076],db_even.mem_bank[2076],db_odd.mem_bank[2077],db_even.mem_bank[2077],db_odd.mem_bank[2078],db_even.mem_bank[2078],db_odd.mem_bank[2079],db_even.mem_bank[2079],db_odd.mem_bank[2080],db_even.mem_bank[2080],db_odd.mem_bank[2081],db_even.mem_bank[2081],db_odd.mem_bank[2082],db_even.mem_bank[2082],db_odd.mem_bank[2083],db_even.mem_bank[2083],db_odd.mem_bank[2084],db_even.mem_bank[2084],db_odd.mem_bank[2085],db_even.mem_bank[2085],db_odd.mem_bank[2086],db_even.mem_bank[2086],db_odd.mem_bank[2087],db_even.mem_bank[2087],db_odd.mem_bank[2088],db_even.mem_bank[2088],db_odd.mem_bank[2089],db_even.mem_bank[2089],db_odd.mem_bank[2090],db_even.mem_bank[2090],db_odd.mem_bank[2091],db_even.mem_bank[2091],db_odd.mem_bank[2092],db_even.mem_bank[2092],db_odd.mem_bank[2093],db_even.mem_bank[2093],db_odd.mem_bank[2094],db_even.mem_bank[2094],db_odd.mem_bank[2095],db_even.mem_bank[2095],db_odd.mem_bank[2096],db_even.mem_bank[2096],db_odd.mem_bank[2097],db_even.mem_bank[2097],db_odd.mem_bank[2098],db_even.mem_bank[2098],db_odd.mem_bank[2099],db_even.mem_bank[2099],db_odd.mem_bank[2100],db_even.mem_bank[2100],db_odd.mem_bank[2101],db_even.mem_bank[2101],db_odd.mem_bank[2102],db_even.mem_bank[2102],db_odd.mem_bank[2103],db_even.mem_bank[2103],db_odd.mem_bank[2104],db_even.mem_bank[2104],db_odd.mem_bank[2105],db_even.mem_bank[2105],db_odd.mem_bank[2106],db_even.mem_bank[2106],db_odd.mem_bank[2107],db_even.mem_bank[2107],db_odd.mem_bank[2108],db_even.mem_bank[2108],db_odd.mem_bank[2109],db_even.mem_bank[2109],db_odd.mem_bank[2110],db_even.mem_bank[2110],db_odd.mem_bank[2111],db_even.mem_bank[2111],db_odd.mem_bank[2112],db_even.mem_bank[2112],db_odd.mem_bank[2113],db_even.mem_bank[2113],db_odd.mem_bank[2114],db_even.mem_bank[2114],db_odd.mem_bank[2115],db_even.mem_bank[2115],db_odd.mem_bank[2116],db_even.mem_bank[2116],db_odd.mem_bank[2117],db_even.mem_bank[2117],db_odd.mem_bank[2118],db_even.mem_bank[2118],db_odd.mem_bank[2119],db_even.mem_bank[2119],db_odd.mem_bank[2120],db_even.mem_bank[2120],db_odd.mem_bank[2121],db_even.mem_bank[2121],db_odd.mem_bank[2122],db_even.mem_bank[2122],db_odd.mem_bank[2123],db_even.mem_bank[2123],db_odd.mem_bank[2124],db_even.mem_bank[2124],db_odd.mem_bank[2125],db_even.mem_bank[2125],db_odd.mem_bank[2126],db_even.mem_bank[2126],db_odd.mem_bank[2127],db_even.mem_bank[2127],db_odd.mem_bank[2128],db_even.mem_bank[2128],db_odd.mem_bank[2129],db_even.mem_bank[2129],db_odd.mem_bank[2130],db_even.mem_bank[2130],db_odd.mem_bank[2131],db_even.mem_bank[2131],db_odd.mem_bank[2132],db_even.mem_bank[2132],db_odd.mem_bank[2133],db_even.mem_bank[2133],db_odd.mem_bank[2134],db_even.mem_bank[2134],db_odd.mem_bank[2135],db_even.mem_bank[2135],db_odd.mem_bank[2136],db_even.mem_bank[2136],db_odd.mem_bank[2137],db_even.mem_bank[2137],db_odd.mem_bank[2138],db_even.mem_bank[2138],db_odd.mem_bank[2139],db_even.mem_bank[2139],db_odd.mem_bank[2140],db_even.mem_bank[2140],db_odd.mem_bank[2141],db_even.mem_bank[2141],db_odd.mem_bank[2142],db_even.mem_bank[2142],db_odd.mem_bank[2143],db_even.mem_bank[2143],db_odd.mem_bank[2144],db_even.mem_bank[2144],db_odd.mem_bank[2145],db_even.mem_bank[2145],db_odd.mem_bank[2146],db_even.mem_bank[2146],db_odd.mem_bank[2147],db_even.mem_bank[2147],db_odd.mem_bank[2148],db_even.mem_bank[2148],db_odd.mem_bank[2149],db_even.mem_bank[2149],db_odd.mem_bank[2150],db_even.mem_bank[2150],db_odd.mem_bank[2151],db_even.mem_bank[2151],db_odd.mem_bank[2152],db_even.mem_bank[2152],db_odd.mem_bank[2153],db_even.mem_bank[2153],db_odd.mem_bank[2154],db_even.mem_bank[2154],db_odd.mem_bank[2155],db_even.mem_bank[2155],db_odd.mem_bank[2156],db_even.mem_bank[2156],db_odd.mem_bank[2157],db_even.mem_bank[2157],db_odd.mem_bank[2158],db_even.mem_bank[2158],db_odd.mem_bank[2159],db_even.mem_bank[2159],db_odd.mem_bank[2160],db_even.mem_bank[2160],db_odd.mem_bank[2161],db_even.mem_bank[2161],db_odd.mem_bank[2162],db_even.mem_bank[2162],db_odd.mem_bank[2163],db_even.mem_bank[2163],db_odd.mem_bank[2164],db_even.mem_bank[2164],db_odd.mem_bank[2165],db_even.mem_bank[2165],db_odd.mem_bank[2166],db_even.mem_bank[2166],db_odd.mem_bank[2167],db_even.mem_bank[2167],db_odd.mem_bank[2168],db_even.mem_bank[2168],db_odd.mem_bank[2169],db_even.mem_bank[2169],db_odd.mem_bank[2170],db_even.mem_bank[2170],db_odd.mem_bank[2171],db_even.mem_bank[2171],db_odd.mem_bank[2172],db_even.mem_bank[2172],db_odd.mem_bank[2173],db_even.mem_bank[2173],db_odd.mem_bank[2174],db_even.mem_bank[2174],db_odd.mem_bank[2175],db_even.mem_bank[2175],db_odd.mem_bank[2176],db_even.mem_bank[2176],db_odd.mem_bank[2177],db_even.mem_bank[2177],db_odd.mem_bank[2178],db_even.mem_bank[2178],db_odd.mem_bank[2179],db_even.mem_bank[2179],db_odd.mem_bank[2180],db_even.mem_bank[2180],db_odd.mem_bank[2181],db_even.mem_bank[2181],db_odd.mem_bank[2182],db_even.mem_bank[2182],db_odd.mem_bank[2183],db_even.mem_bank[2183],db_odd.mem_bank[2184],db_even.mem_bank[2184],db_odd.mem_bank[2185],db_even.mem_bank[2185],db_odd.mem_bank[2186],db_even.mem_bank[2186],db_odd.mem_bank[2187],db_even.mem_bank[2187],db_odd.mem_bank[2188],db_even.mem_bank[2188],db_odd.mem_bank[2189],db_even.mem_bank[2189],db_odd.mem_bank[2190],db_even.mem_bank[2190],db_odd.mem_bank[2191],db_even.mem_bank[2191],db_odd.mem_bank[2192],db_even.mem_bank[2192],db_odd.mem_bank[2193],db_even.mem_bank[2193],db_odd.mem_bank[2194],db_even.mem_bank[2194],db_odd.mem_bank[2195],db_even.mem_bank[2195],db_odd.mem_bank[2196],db_even.mem_bank[2196],db_odd.mem_bank[2197],db_even.mem_bank[2197],db_odd.mem_bank[2198],db_even.mem_bank[2198],db_odd.mem_bank[2199],db_even.mem_bank[2199],db_odd.mem_bank[2200],db_even.mem_bank[2200],db_odd.mem_bank[2201],db_even.mem_bank[2201],db_odd.mem_bank[2202],db_even.mem_bank[2202],db_odd.mem_bank[2203],db_even.mem_bank[2203],db_odd.mem_bank[2204],db_even.mem_bank[2204],db_odd.mem_bank[2205],db_even.mem_bank[2205],db_odd.mem_bank[2206],db_even.mem_bank[2206],db_odd.mem_bank[2207],db_even.mem_bank[2207],db_odd.mem_bank[2208],db_even.mem_bank[2208],db_odd.mem_bank[2209],db_even.mem_bank[2209],db_odd.mem_bank[2210],db_even.mem_bank[2210],db_odd.mem_bank[2211],db_even.mem_bank[2211],db_odd.mem_bank[2212],db_even.mem_bank[2212],db_odd.mem_bank[2213],db_even.mem_bank[2213],db_odd.mem_bank[2214],db_even.mem_bank[2214],db_odd.mem_bank[2215],db_even.mem_bank[2215],db_odd.mem_bank[2216],db_even.mem_bank[2216],db_odd.mem_bank[2217],db_even.mem_bank[2217],db_odd.mem_bank[2218],db_even.mem_bank[2218],db_odd.mem_bank[2219],db_even.mem_bank[2219],db_odd.mem_bank[2220],db_even.mem_bank[2220],db_odd.mem_bank[2221],db_even.mem_bank[2221],db_odd.mem_bank[2222],db_even.mem_bank[2222],db_odd.mem_bank[2223],db_even.mem_bank[2223],db_odd.mem_bank[2224],db_even.mem_bank[2224],db_odd.mem_bank[2225],db_even.mem_bank[2225],db_odd.mem_bank[2226],db_even.mem_bank[2226],db_odd.mem_bank[2227],db_even.mem_bank[2227],db_odd.mem_bank[2228],db_even.mem_bank[2228],db_odd.mem_bank[2229],db_even.mem_bank[2229],db_odd.mem_bank[2230],db_even.mem_bank[2230],db_odd.mem_bank[2231],db_even.mem_bank[2231],db_odd.mem_bank[2232],db_even.mem_bank[2232],db_odd.mem_bank[2233],db_even.mem_bank[2233],db_odd.mem_bank[2234],db_even.mem_bank[2234],db_odd.mem_bank[2235],db_even.mem_bank[2235],db_odd.mem_bank[2236],db_even.mem_bank[2236],db_odd.mem_bank[2237],db_even.mem_bank[2237],db_odd.mem_bank[2238],db_even.mem_bank[2238],db_odd.mem_bank[2239],db_even.mem_bank[2239],db_odd.mem_bank[2240],db_even.mem_bank[2240],db_odd.mem_bank[2241],db_even.mem_bank[2241],db_odd.mem_bank[2242],db_even.mem_bank[2242],db_odd.mem_bank[2243],db_even.mem_bank[2243],db_odd.mem_bank[2244],db_even.mem_bank[2244],db_odd.mem_bank[2245],db_even.mem_bank[2245],db_odd.mem_bank[2246],db_even.mem_bank[2246],db_odd.mem_bank[2247],db_even.mem_bank[2247],db_odd.mem_bank[2248],db_even.mem_bank[2248],db_odd.mem_bank[2249],db_even.mem_bank[2249],db_odd.mem_bank[2250],db_even.mem_bank[2250],db_odd.mem_bank[2251],db_even.mem_bank[2251],db_odd.mem_bank[2252],db_even.mem_bank[2252],db_odd.mem_bank[2253],db_even.mem_bank[2253],db_odd.mem_bank[2254],db_even.mem_bank[2254],db_odd.mem_bank[2255],db_even.mem_bank[2255],db_odd.mem_bank[2256],db_even.mem_bank[2256],db_odd.mem_bank[2257],db_even.mem_bank[2257],db_odd.mem_bank[2258],db_even.mem_bank[2258],db_odd.mem_bank[2259],db_even.mem_bank[2259],db_odd.mem_bank[2260],db_even.mem_bank[2260],db_odd.mem_bank[2261],db_even.mem_bank[2261],db_odd.mem_bank[2262],db_even.mem_bank[2262],db_odd.mem_bank[2263],db_even.mem_bank[2263],db_odd.mem_bank[2264],db_even.mem_bank[2264],db_odd.mem_bank[2265],db_even.mem_bank[2265],db_odd.mem_bank[2266],db_even.mem_bank[2266],db_odd.mem_bank[2267],db_even.mem_bank[2267],db_odd.mem_bank[2268],db_even.mem_bank[2268],db_odd.mem_bank[2269],db_even.mem_bank[2269],db_odd.mem_bank[2270],db_even.mem_bank[2270],db_odd.mem_bank[2271],db_even.mem_bank[2271],db_odd.mem_bank[2272],db_even.mem_bank[2272],db_odd.mem_bank[2273],db_even.mem_bank[2273],db_odd.mem_bank[2274],db_even.mem_bank[2274],db_odd.mem_bank[2275],db_even.mem_bank[2275],db_odd.mem_bank[2276],db_even.mem_bank[2276],db_odd.mem_bank[2277],db_even.mem_bank[2277],db_odd.mem_bank[2278],db_even.mem_bank[2278],db_odd.mem_bank[2279],db_even.mem_bank[2279],db_odd.mem_bank[2280],db_even.mem_bank[2280],db_odd.mem_bank[2281],db_even.mem_bank[2281],db_odd.mem_bank[2282],db_even.mem_bank[2282],db_odd.mem_bank[2283],db_even.mem_bank[2283],db_odd.mem_bank[2284],db_even.mem_bank[2284],db_odd.mem_bank[2285],db_even.mem_bank[2285],db_odd.mem_bank[2286],db_even.mem_bank[2286],db_odd.mem_bank[2287],db_even.mem_bank[2287],db_odd.mem_bank[2288],db_even.mem_bank[2288],db_odd.mem_bank[2289],db_even.mem_bank[2289],db_odd.mem_bank[2290],db_even.mem_bank[2290],db_odd.mem_bank[2291],db_even.mem_bank[2291],db_odd.mem_bank[2292],db_even.mem_bank[2292],db_odd.mem_bank[2293],db_even.mem_bank[2293],db_odd.mem_bank[2294],db_even.mem_bank[2294],db_odd.mem_bank[2295],db_even.mem_bank[2295],db_odd.mem_bank[2296],db_even.mem_bank[2296],db_odd.mem_bank[2297],db_even.mem_bank[2297],db_odd.mem_bank[2298],db_even.mem_bank[2298],db_odd.mem_bank[2299],db_even.mem_bank[2299],db_odd.mem_bank[2300],db_even.mem_bank[2300],db_odd.mem_bank[2301],db_even.mem_bank[2301],db_odd.mem_bank[2302],db_even.mem_bank[2302],db_odd.mem_bank[2303],db_even.mem_bank[2303],db_odd.mem_bank[2304],db_even.mem_bank[2304],db_odd.mem_bank[2305],db_even.mem_bank[2305],db_odd.mem_bank[2306],db_even.mem_bank[2306],db_odd.mem_bank[2307],db_even.mem_bank[2307],db_odd.mem_bank[2308],db_even.mem_bank[2308],db_odd.mem_bank[2309],db_even.mem_bank[2309],db_odd.mem_bank[2310],db_even.mem_bank[2310],db_odd.mem_bank[2311],db_even.mem_bank[2311],db_odd.mem_bank[2312],db_even.mem_bank[2312],db_odd.mem_bank[2313],db_even.mem_bank[2313],db_odd.mem_bank[2314],db_even.mem_bank[2314],db_odd.mem_bank[2315],db_even.mem_bank[2315],db_odd.mem_bank[2316],db_even.mem_bank[2316],db_odd.mem_bank[2317],db_even.mem_bank[2317],db_odd.mem_bank[2318],db_even.mem_bank[2318],db_odd.mem_bank[2319],db_even.mem_bank[2319],db_odd.mem_bank[2320],db_even.mem_bank[2320],db_odd.mem_bank[2321],db_even.mem_bank[2321],db_odd.mem_bank[2322],db_even.mem_bank[2322],db_odd.mem_bank[2323],db_even.mem_bank[2323],db_odd.mem_bank[2324],db_even.mem_bank[2324],db_odd.mem_bank[2325],db_even.mem_bank[2325],db_odd.mem_bank[2326],db_even.mem_bank[2326],db_odd.mem_bank[2327],db_even.mem_bank[2327],db_odd.mem_bank[2328],db_even.mem_bank[2328],db_odd.mem_bank[2329],db_even.mem_bank[2329],db_odd.mem_bank[2330],db_even.mem_bank[2330],db_odd.mem_bank[2331],db_even.mem_bank[2331],db_odd.mem_bank[2332],db_even.mem_bank[2332],db_odd.mem_bank[2333],db_even.mem_bank[2333],db_odd.mem_bank[2334],db_even.mem_bank[2334],db_odd.mem_bank[2335],db_even.mem_bank[2335],db_odd.mem_bank[2336],db_even.mem_bank[2336],db_odd.mem_bank[2337],db_even.mem_bank[2337],db_odd.mem_bank[2338],db_even.mem_bank[2338],db_odd.mem_bank[2339],db_even.mem_bank[2339],db_odd.mem_bank[2340],db_even.mem_bank[2340],db_odd.mem_bank[2341],db_even.mem_bank[2341],db_odd.mem_bank[2342],db_even.mem_bank[2342],db_odd.mem_bank[2343],db_even.mem_bank[2343],db_odd.mem_bank[2344],db_even.mem_bank[2344],db_odd.mem_bank[2345],db_even.mem_bank[2345],db_odd.mem_bank[2346],db_even.mem_bank[2346],db_odd.mem_bank[2347],db_even.mem_bank[2347],db_odd.mem_bank[2348],db_even.mem_bank[2348],db_odd.mem_bank[2349],db_even.mem_bank[2349],db_odd.mem_bank[2350],db_even.mem_bank[2350],db_odd.mem_bank[2351],db_even.mem_bank[2351],db_odd.mem_bank[2352],db_even.mem_bank[2352],db_odd.mem_bank[2353],db_even.mem_bank[2353],db_odd.mem_bank[2354],db_even.mem_bank[2354],db_odd.mem_bank[2355],db_even.mem_bank[2355],db_odd.mem_bank[2356],db_even.mem_bank[2356],db_odd.mem_bank[2357],db_even.mem_bank[2357],db_odd.mem_bank[2358],db_even.mem_bank[2358],db_odd.mem_bank[2359],db_even.mem_bank[2359],db_odd.mem_bank[2360],db_even.mem_bank[2360],db_odd.mem_bank[2361],db_even.mem_bank[2361],db_odd.mem_bank[2362],db_even.mem_bank[2362],db_odd.mem_bank[2363],db_even.mem_bank[2363],db_odd.mem_bank[2364],db_even.mem_bank[2364],db_odd.mem_bank[2365],db_even.mem_bank[2365],db_odd.mem_bank[2366],db_even.mem_bank[2366],db_odd.mem_bank[2367],db_even.mem_bank[2367],db_odd.mem_bank[2368],db_even.mem_bank[2368],db_odd.mem_bank[2369],db_even.mem_bank[2369],db_odd.mem_bank[2370],db_even.mem_bank[2370],db_odd.mem_bank[2371],db_even.mem_bank[2371],db_odd.mem_bank[2372],db_even.mem_bank[2372],db_odd.mem_bank[2373],db_even.mem_bank[2373],db_odd.mem_bank[2374],db_even.mem_bank[2374],db_odd.mem_bank[2375],db_even.mem_bank[2375],db_odd.mem_bank[2376],db_even.mem_bank[2376],db_odd.mem_bank[2377],db_even.mem_bank[2377],db_odd.mem_bank[2378],db_even.mem_bank[2378],db_odd.mem_bank[2379],db_even.mem_bank[2379],db_odd.mem_bank[2380],db_even.mem_bank[2380],db_odd.mem_bank[2381],db_even.mem_bank[2381],db_odd.mem_bank[2382],db_even.mem_bank[2382],db_odd.mem_bank[2383],db_even.mem_bank[2383],db_odd.mem_bank[2384],db_even.mem_bank[2384],db_odd.mem_bank[2385],db_even.mem_bank[2385],db_odd.mem_bank[2386],db_even.mem_bank[2386],db_odd.mem_bank[2387],db_even.mem_bank[2387],db_odd.mem_bank[2388],db_even.mem_bank[2388],db_odd.mem_bank[2389],db_even.mem_bank[2389],db_odd.mem_bank[2390],db_even.mem_bank[2390],db_odd.mem_bank[2391],db_even.mem_bank[2391],db_odd.mem_bank[2392],db_even.mem_bank[2392],db_odd.mem_bank[2393],db_even.mem_bank[2393],db_odd.mem_bank[2394],db_even.mem_bank[2394],db_odd.mem_bank[2395],db_even.mem_bank[2395],db_odd.mem_bank[2396],db_even.mem_bank[2396],db_odd.mem_bank[2397],db_even.mem_bank[2397],db_odd.mem_bank[2398],db_even.mem_bank[2398],db_odd.mem_bank[2399],db_even.mem_bank[2399],db_odd.mem_bank[2400],db_even.mem_bank[2400],db_odd.mem_bank[2401],db_even.mem_bank[2401],db_odd.mem_bank[2402],db_even.mem_bank[2402],db_odd.mem_bank[2403],db_even.mem_bank[2403],db_odd.mem_bank[2404],db_even.mem_bank[2404],db_odd.mem_bank[2405],db_even.mem_bank[2405],db_odd.mem_bank[2406],db_even.mem_bank[2406],db_odd.mem_bank[2407],db_even.mem_bank[2407],db_odd.mem_bank[2408],db_even.mem_bank[2408],db_odd.mem_bank[2409],db_even.mem_bank[2409],db_odd.mem_bank[2410],db_even.mem_bank[2410],db_odd.mem_bank[2411],db_even.mem_bank[2411],db_odd.mem_bank[2412],db_even.mem_bank[2412],db_odd.mem_bank[2413],db_even.mem_bank[2413],db_odd.mem_bank[2414],db_even.mem_bank[2414],db_odd.mem_bank[2415],db_even.mem_bank[2415],db_odd.mem_bank[2416],db_even.mem_bank[2416],db_odd.mem_bank[2417],db_even.mem_bank[2417],db_odd.mem_bank[2418],db_even.mem_bank[2418],db_odd.mem_bank[2419],db_even.mem_bank[2419],db_odd.mem_bank[2420],db_even.mem_bank[2420],db_odd.mem_bank[2421],db_even.mem_bank[2421],db_odd.mem_bank[2422],db_even.mem_bank[2422],db_odd.mem_bank[2423],db_even.mem_bank[2423],db_odd.mem_bank[2424],db_even.mem_bank[2424],db_odd.mem_bank[2425],db_even.mem_bank[2425],db_odd.mem_bank[2426],db_even.mem_bank[2426],db_odd.mem_bank[2427],db_even.mem_bank[2427],db_odd.mem_bank[2428],db_even.mem_bank[2428],db_odd.mem_bank[2429],db_even.mem_bank[2429],db_odd.mem_bank[2430],db_even.mem_bank[2430],db_odd.mem_bank[2431],db_even.mem_bank[2431],db_odd.mem_bank[2432],db_even.mem_bank[2432],db_odd.mem_bank[2433],db_even.mem_bank[2433],db_odd.mem_bank[2434],db_even.mem_bank[2434],db_odd.mem_bank[2435],db_even.mem_bank[2435],db_odd.mem_bank[2436],db_even.mem_bank[2436],db_odd.mem_bank[2437],db_even.mem_bank[2437],db_odd.mem_bank[2438],db_even.mem_bank[2438],db_odd.mem_bank[2439],db_even.mem_bank[2439],db_odd.mem_bank[2440],db_even.mem_bank[2440],db_odd.mem_bank[2441],db_even.mem_bank[2441],db_odd.mem_bank[2442],db_even.mem_bank[2442],db_odd.mem_bank[2443],db_even.mem_bank[2443],db_odd.mem_bank[2444],db_even.mem_bank[2444],db_odd.mem_bank[2445],db_even.mem_bank[2445],db_odd.mem_bank[2446],db_even.mem_bank[2446],db_odd.mem_bank[2447],db_even.mem_bank[2447],db_odd.mem_bank[2448],db_even.mem_bank[2448],db_odd.mem_bank[2449],db_even.mem_bank[2449],db_odd.mem_bank[2450],db_even.mem_bank[2450],db_odd.mem_bank[2451],db_even.mem_bank[2451],db_odd.mem_bank[2452],db_even.mem_bank[2452],db_odd.mem_bank[2453],db_even.mem_bank[2453],db_odd.mem_bank[2454],db_even.mem_bank[2454],db_odd.mem_bank[2455],db_even.mem_bank[2455],db_odd.mem_bank[2456],db_even.mem_bank[2456],db_odd.mem_bank[2457],db_even.mem_bank[2457],db_odd.mem_bank[2458],db_even.mem_bank[2458],db_odd.mem_bank[2459],db_even.mem_bank[2459],db_odd.mem_bank[2460],db_even.mem_bank[2460],db_odd.mem_bank[2461],db_even.mem_bank[2461],db_odd.mem_bank[2462],db_even.mem_bank[2462],db_odd.mem_bank[2463],db_even.mem_bank[2463],db_odd.mem_bank[2464],db_even.mem_bank[2464],db_odd.mem_bank[2465],db_even.mem_bank[2465],db_odd.mem_bank[2466],db_even.mem_bank[2466],db_odd.mem_bank[2467],db_even.mem_bank[2467],db_odd.mem_bank[2468],db_even.mem_bank[2468],db_odd.mem_bank[2469],db_even.mem_bank[2469],db_odd.mem_bank[2470],db_even.mem_bank[2470],db_odd.mem_bank[2471],db_even.mem_bank[2471],db_odd.mem_bank[2472],db_even.mem_bank[2472],db_odd.mem_bank[2473],db_even.mem_bank[2473],db_odd.mem_bank[2474],db_even.mem_bank[2474],db_odd.mem_bank[2475],db_even.mem_bank[2475],db_odd.mem_bank[2476],db_even.mem_bank[2476],db_odd.mem_bank[2477],db_even.mem_bank[2477],db_odd.mem_bank[2478],db_even.mem_bank[2478],db_odd.mem_bank[2479],db_even.mem_bank[2479],db_odd.mem_bank[2480],db_even.mem_bank[2480],db_odd.mem_bank[2481],db_even.mem_bank[2481],db_odd.mem_bank[2482],db_even.mem_bank[2482],db_odd.mem_bank[2483],db_even.mem_bank[2483],db_odd.mem_bank[2484],db_even.mem_bank[2484],db_odd.mem_bank[2485],db_even.mem_bank[2485],db_odd.mem_bank[2486],db_even.mem_bank[2486],db_odd.mem_bank[2487],db_even.mem_bank[2487],db_odd.mem_bank[2488],db_even.mem_bank[2488],db_odd.mem_bank[2489],db_even.mem_bank[2489],db_odd.mem_bank[2490],db_even.mem_bank[2490],db_odd.mem_bank[2491],db_even.mem_bank[2491],db_odd.mem_bank[2492],db_even.mem_bank[2492],db_odd.mem_bank[2493],db_even.mem_bank[2493],db_odd.mem_bank[2494],db_even.mem_bank[2494],db_odd.mem_bank[2495],db_even.mem_bank[2495],db_odd.mem_bank[2496],db_even.mem_bank[2496],db_odd.mem_bank[2497],db_even.mem_bank[2497],db_odd.mem_bank[2498],db_even.mem_bank[2498],db_odd.mem_bank[2499],db_even.mem_bank[2499],db_odd.mem_bank[2500],db_even.mem_bank[2500],db_odd.mem_bank[2501],db_even.mem_bank[2501],db_odd.mem_bank[2502],db_even.mem_bank[2502],db_odd.mem_bank[2503],db_even.mem_bank[2503],db_odd.mem_bank[2504],db_even.mem_bank[2504],db_odd.mem_bank[2505],db_even.mem_bank[2505],db_odd.mem_bank[2506],db_even.mem_bank[2506],db_odd.mem_bank[2507],db_even.mem_bank[2507],db_odd.mem_bank[2508],db_even.mem_bank[2508],db_odd.mem_bank[2509],db_even.mem_bank[2509],db_odd.mem_bank[2510],db_even.mem_bank[2510],db_odd.mem_bank[2511],db_even.mem_bank[2511],db_odd.mem_bank[2512],db_even.mem_bank[2512],db_odd.mem_bank[2513],db_even.mem_bank[2513],db_odd.mem_bank[2514],db_even.mem_bank[2514],db_odd.mem_bank[2515],db_even.mem_bank[2515],db_odd.mem_bank[2516],db_even.mem_bank[2516],db_odd.mem_bank[2517],db_even.mem_bank[2517],db_odd.mem_bank[2518],db_even.mem_bank[2518],db_odd.mem_bank[2519],db_even.mem_bank[2519],db_odd.mem_bank[2520],db_even.mem_bank[2520],db_odd.mem_bank[2521],db_even.mem_bank[2521],db_odd.mem_bank[2522],db_even.mem_bank[2522],db_odd.mem_bank[2523],db_even.mem_bank[2523],db_odd.mem_bank[2524],db_even.mem_bank[2524],db_odd.mem_bank[2525],db_even.mem_bank[2525],db_odd.mem_bank[2526],db_even.mem_bank[2526],db_odd.mem_bank[2527],db_even.mem_bank[2527],db_odd.mem_bank[2528],db_even.mem_bank[2528],db_odd.mem_bank[2529],db_even.mem_bank[2529],db_odd.mem_bank[2530],db_even.mem_bank[2530],db_odd.mem_bank[2531],db_even.mem_bank[2531],db_odd.mem_bank[2532],db_even.mem_bank[2532],db_odd.mem_bank[2533],db_even.mem_bank[2533],db_odd.mem_bank[2534],db_even.mem_bank[2534],db_odd.mem_bank[2535],db_even.mem_bank[2535],db_odd.mem_bank[2536],db_even.mem_bank[2536],db_odd.mem_bank[2537],db_even.mem_bank[2537],db_odd.mem_bank[2538],db_even.mem_bank[2538],db_odd.mem_bank[2539],db_even.mem_bank[2539],db_odd.mem_bank[2540],db_even.mem_bank[2540],db_odd.mem_bank[2541],db_even.mem_bank[2541],db_odd.mem_bank[2542],db_even.mem_bank[2542],db_odd.mem_bank[2543],db_even.mem_bank[2543],db_odd.mem_bank[2544],db_even.mem_bank[2544],db_odd.mem_bank[2545],db_even.mem_bank[2545],db_odd.mem_bank[2546],db_even.mem_bank[2546],db_odd.mem_bank[2547],db_even.mem_bank[2547],db_odd.mem_bank[2548],db_even.mem_bank[2548],db_odd.mem_bank[2549],db_even.mem_bank[2549],db_odd.mem_bank[2550],db_even.mem_bank[2550],db_odd.mem_bank[2551],db_even.mem_bank[2551],db_odd.mem_bank[2552],db_even.mem_bank[2552],db_odd.mem_bank[2553],db_even.mem_bank[2553],db_odd.mem_bank[2554],db_even.mem_bank[2554],db_odd.mem_bank[2555],db_even.mem_bank[2555],db_odd.mem_bank[2556],db_even.mem_bank[2556],db_odd.mem_bank[2557],db_even.mem_bank[2557],db_odd.mem_bank[2558],db_even.mem_bank[2558],db_odd.mem_bank[2559],db_even.mem_bank[2559],db_odd.mem_bank[2560],db_even.mem_bank[2560],db_odd.mem_bank[2561],db_even.mem_bank[2561],db_odd.mem_bank[2562],db_even.mem_bank[2562],db_odd.mem_bank[2563],db_even.mem_bank[2563],db_odd.mem_bank[2564],db_even.mem_bank[2564],db_odd.mem_bank[2565],db_even.mem_bank[2565],db_odd.mem_bank[2566],db_even.mem_bank[2566],db_odd.mem_bank[2567],db_even.mem_bank[2567],db_odd.mem_bank[2568],db_even.mem_bank[2568],db_odd.mem_bank[2569],db_even.mem_bank[2569],db_odd.mem_bank[2570],db_even.mem_bank[2570],db_odd.mem_bank[2571],db_even.mem_bank[2571],db_odd.mem_bank[2572],db_even.mem_bank[2572],db_odd.mem_bank[2573],db_even.mem_bank[2573],db_odd.mem_bank[2574],db_even.mem_bank[2574],db_odd.mem_bank[2575],db_even.mem_bank[2575],db_odd.mem_bank[2576],db_even.mem_bank[2576],db_odd.mem_bank[2577],db_even.mem_bank[2577],db_odd.mem_bank[2578],db_even.mem_bank[2578],db_odd.mem_bank[2579],db_even.mem_bank[2579],db_odd.mem_bank[2580],db_even.mem_bank[2580],db_odd.mem_bank[2581],db_even.mem_bank[2581],db_odd.mem_bank[2582],db_even.mem_bank[2582],db_odd.mem_bank[2583],db_even.mem_bank[2583],db_odd.mem_bank[2584],db_even.mem_bank[2584],db_odd.mem_bank[2585],db_even.mem_bank[2585],db_odd.mem_bank[2586],db_even.mem_bank[2586],db_odd.mem_bank[2587],db_even.mem_bank[2587],db_odd.mem_bank[2588],db_even.mem_bank[2588],db_odd.mem_bank[2589],db_even.mem_bank[2589],db_odd.mem_bank[2590],db_even.mem_bank[2590],db_odd.mem_bank[2591],db_even.mem_bank[2591],db_odd.mem_bank[2592],db_even.mem_bank[2592],db_odd.mem_bank[2593],db_even.mem_bank[2593],db_odd.mem_bank[2594],db_even.mem_bank[2594],db_odd.mem_bank[2595],db_even.mem_bank[2595],db_odd.mem_bank[2596],db_even.mem_bank[2596],db_odd.mem_bank[2597],db_even.mem_bank[2597],db_odd.mem_bank[2598],db_even.mem_bank[2598],db_odd.mem_bank[2599],db_even.mem_bank[2599],db_odd.mem_bank[2600],db_even.mem_bank[2600],db_odd.mem_bank[2601],db_even.mem_bank[2601],db_odd.mem_bank[2602],db_even.mem_bank[2602],db_odd.mem_bank[2603],db_even.mem_bank[2603],db_odd.mem_bank[2604],db_even.mem_bank[2604],db_odd.mem_bank[2605],db_even.mem_bank[2605],db_odd.mem_bank[2606],db_even.mem_bank[2606],db_odd.mem_bank[2607],db_even.mem_bank[2607],db_odd.mem_bank[2608],db_even.mem_bank[2608],db_odd.mem_bank[2609],db_even.mem_bank[2609],db_odd.mem_bank[2610],db_even.mem_bank[2610],db_odd.mem_bank[2611],db_even.mem_bank[2611],db_odd.mem_bank[2612],db_even.mem_bank[2612],db_odd.mem_bank[2613],db_even.mem_bank[2613],db_odd.mem_bank[2614],db_even.mem_bank[2614],db_odd.mem_bank[2615],db_even.mem_bank[2615],db_odd.mem_bank[2616],db_even.mem_bank[2616],db_odd.mem_bank[2617],db_even.mem_bank[2617],db_odd.mem_bank[2618],db_even.mem_bank[2618],db_odd.mem_bank[2619],db_even.mem_bank[2619],db_odd.mem_bank[2620],db_even.mem_bank[2620],db_odd.mem_bank[2621],db_even.mem_bank[2621],db_odd.mem_bank[2622],db_even.mem_bank[2622],db_odd.mem_bank[2623],db_even.mem_bank[2623],db_odd.mem_bank[2624],db_even.mem_bank[2624],db_odd.mem_bank[2625],db_even.mem_bank[2625],db_odd.mem_bank[2626],db_even.mem_bank[2626],db_odd.mem_bank[2627],db_even.mem_bank[2627],db_odd.mem_bank[2628],db_even.mem_bank[2628],db_odd.mem_bank[2629],db_even.mem_bank[2629],db_odd.mem_bank[2630],db_even.mem_bank[2630],db_odd.mem_bank[2631],db_even.mem_bank[2631],db_odd.mem_bank[2632],db_even.mem_bank[2632],db_odd.mem_bank[2633],db_even.mem_bank[2633],db_odd.mem_bank[2634],db_even.mem_bank[2634],db_odd.mem_bank[2635],db_even.mem_bank[2635],db_odd.mem_bank[2636],db_even.mem_bank[2636],db_odd.mem_bank[2637],db_even.mem_bank[2637],db_odd.mem_bank[2638],db_even.mem_bank[2638],db_odd.mem_bank[2639],db_even.mem_bank[2639],db_odd.mem_bank[2640],db_even.mem_bank[2640],db_odd.mem_bank[2641],db_even.mem_bank[2641],db_odd.mem_bank[2642],db_even.mem_bank[2642],db_odd.mem_bank[2643],db_even.mem_bank[2643],db_odd.mem_bank[2644],db_even.mem_bank[2644],db_odd.mem_bank[2645],db_even.mem_bank[2645],db_odd.mem_bank[2646],db_even.mem_bank[2646],db_odd.mem_bank[2647],db_even.mem_bank[2647],db_odd.mem_bank[2648],db_even.mem_bank[2648],db_odd.mem_bank[2649],db_even.mem_bank[2649],db_odd.mem_bank[2650],db_even.mem_bank[2650],db_odd.mem_bank[2651],db_even.mem_bank[2651],db_odd.mem_bank[2652],db_even.mem_bank[2652],db_odd.mem_bank[2653],db_even.mem_bank[2653],db_odd.mem_bank[2654],db_even.mem_bank[2654],db_odd.mem_bank[2655],db_even.mem_bank[2655],db_odd.mem_bank[2656],db_even.mem_bank[2656],db_odd.mem_bank[2657],db_even.mem_bank[2657],db_odd.mem_bank[2658],db_even.mem_bank[2658],db_odd.mem_bank[2659],db_even.mem_bank[2659],db_odd.mem_bank[2660],db_even.mem_bank[2660],db_odd.mem_bank[2661],db_even.mem_bank[2661],db_odd.mem_bank[2662],db_even.mem_bank[2662],db_odd.mem_bank[2663],db_even.mem_bank[2663],db_odd.mem_bank[2664],db_even.mem_bank[2664],db_odd.mem_bank[2665],db_even.mem_bank[2665],db_odd.mem_bank[2666],db_even.mem_bank[2666],db_odd.mem_bank[2667],db_even.mem_bank[2667],db_odd.mem_bank[2668],db_even.mem_bank[2668],db_odd.mem_bank[2669],db_even.mem_bank[2669],db_odd.mem_bank[2670],db_even.mem_bank[2670],db_odd.mem_bank[2671],db_even.mem_bank[2671],db_odd.mem_bank[2672],db_even.mem_bank[2672],db_odd.mem_bank[2673],db_even.mem_bank[2673],db_odd.mem_bank[2674],db_even.mem_bank[2674],db_odd.mem_bank[2675],db_even.mem_bank[2675],db_odd.mem_bank[2676],db_even.mem_bank[2676],db_odd.mem_bank[2677],db_even.mem_bank[2677],db_odd.mem_bank[2678],db_even.mem_bank[2678],db_odd.mem_bank[2679],db_even.mem_bank[2679],db_odd.mem_bank[2680],db_even.mem_bank[2680],db_odd.mem_bank[2681],db_even.mem_bank[2681],db_odd.mem_bank[2682],db_even.mem_bank[2682],db_odd.mem_bank[2683],db_even.mem_bank[2683],db_odd.mem_bank[2684],db_even.mem_bank[2684],db_odd.mem_bank[2685],db_even.mem_bank[2685],db_odd.mem_bank[2686],db_even.mem_bank[2686],db_odd.mem_bank[2687],db_even.mem_bank[2687],db_odd.mem_bank[2688],db_even.mem_bank[2688],db_odd.mem_bank[2689],db_even.mem_bank[2689],db_odd.mem_bank[2690],db_even.mem_bank[2690],db_odd.mem_bank[2691],db_even.mem_bank[2691],db_odd.mem_bank[2692],db_even.mem_bank[2692],db_odd.mem_bank[2693],db_even.mem_bank[2693],db_odd.mem_bank[2694],db_even.mem_bank[2694],db_odd.mem_bank[2695],db_even.mem_bank[2695],db_odd.mem_bank[2696],db_even.mem_bank[2696],db_odd.mem_bank[2697],db_even.mem_bank[2697],db_odd.mem_bank[2698],db_even.mem_bank[2698],db_odd.mem_bank[2699],db_even.mem_bank[2699],db_odd.mem_bank[2700],db_even.mem_bank[2700],db_odd.mem_bank[2701],db_even.mem_bank[2701],db_odd.mem_bank[2702],db_even.mem_bank[2702],db_odd.mem_bank[2703],db_even.mem_bank[2703],db_odd.mem_bank[2704],db_even.mem_bank[2704],db_odd.mem_bank[2705],db_even.mem_bank[2705],db_odd.mem_bank[2706],db_even.mem_bank[2706],db_odd.mem_bank[2707],db_even.mem_bank[2707],db_odd.mem_bank[2708],db_even.mem_bank[2708],db_odd.mem_bank[2709],db_even.mem_bank[2709],db_odd.mem_bank[2710],db_even.mem_bank[2710],db_odd.mem_bank[2711],db_even.mem_bank[2711],db_odd.mem_bank[2712],db_even.mem_bank[2712],db_odd.mem_bank[2713],db_even.mem_bank[2713],db_odd.mem_bank[2714],db_even.mem_bank[2714],db_odd.mem_bank[2715],db_even.mem_bank[2715],db_odd.mem_bank[2716],db_even.mem_bank[2716],db_odd.mem_bank[2717],db_even.mem_bank[2717],db_odd.mem_bank[2718],db_even.mem_bank[2718],db_odd.mem_bank[2719],db_even.mem_bank[2719],db_odd.mem_bank[2720],db_even.mem_bank[2720],db_odd.mem_bank[2721],db_even.mem_bank[2721],db_odd.mem_bank[2722],db_even.mem_bank[2722],db_odd.mem_bank[2723],db_even.mem_bank[2723],db_odd.mem_bank[2724],db_even.mem_bank[2724],db_odd.mem_bank[2725],db_even.mem_bank[2725],db_odd.mem_bank[2726],db_even.mem_bank[2726],db_odd.mem_bank[2727],db_even.mem_bank[2727],db_odd.mem_bank[2728],db_even.mem_bank[2728],db_odd.mem_bank[2729],db_even.mem_bank[2729],db_odd.mem_bank[2730],db_even.mem_bank[2730],db_odd.mem_bank[2731],db_even.mem_bank[2731],db_odd.mem_bank[2732],db_even.mem_bank[2732],db_odd.mem_bank[2733],db_even.mem_bank[2733],db_odd.mem_bank[2734],db_even.mem_bank[2734],db_odd.mem_bank[2735],db_even.mem_bank[2735],db_odd.mem_bank[2736],db_even.mem_bank[2736],db_odd.mem_bank[2737],db_even.mem_bank[2737],db_odd.mem_bank[2738],db_even.mem_bank[2738],db_odd.mem_bank[2739],db_even.mem_bank[2739],db_odd.mem_bank[2740],db_even.mem_bank[2740],db_odd.mem_bank[2741],db_even.mem_bank[2741],db_odd.mem_bank[2742],db_even.mem_bank[2742],db_odd.mem_bank[2743],db_even.mem_bank[2743],db_odd.mem_bank[2744],db_even.mem_bank[2744],db_odd.mem_bank[2745],db_even.mem_bank[2745],db_odd.mem_bank[2746],db_even.mem_bank[2746],db_odd.mem_bank[2747],db_even.mem_bank[2747],db_odd.mem_bank[2748],db_even.mem_bank[2748],db_odd.mem_bank[2749],db_even.mem_bank[2749],db_odd.mem_bank[2750],db_even.mem_bank[2750],db_odd.mem_bank[2751],db_even.mem_bank[2751],db_odd.mem_bank[2752],db_even.mem_bank[2752],db_odd.mem_bank[2753],db_even.mem_bank[2753],db_odd.mem_bank[2754],db_even.mem_bank[2754],db_odd.mem_bank[2755],db_even.mem_bank[2755],db_odd.mem_bank[2756],db_even.mem_bank[2756],db_odd.mem_bank[2757],db_even.mem_bank[2757],db_odd.mem_bank[2758],db_even.mem_bank[2758],db_odd.mem_bank[2759],db_even.mem_bank[2759],db_odd.mem_bank[2760],db_even.mem_bank[2760],db_odd.mem_bank[2761],db_even.mem_bank[2761],db_odd.mem_bank[2762],db_even.mem_bank[2762],db_odd.mem_bank[2763],db_even.mem_bank[2763],db_odd.mem_bank[2764],db_even.mem_bank[2764],db_odd.mem_bank[2765],db_even.mem_bank[2765],db_odd.mem_bank[2766],db_even.mem_bank[2766],db_odd.mem_bank[2767],db_even.mem_bank[2767],db_odd.mem_bank[2768],db_even.mem_bank[2768],db_odd.mem_bank[2769],db_even.mem_bank[2769],db_odd.mem_bank[2770],db_even.mem_bank[2770],db_odd.mem_bank[2771],db_even.mem_bank[2771],db_odd.mem_bank[2772],db_even.mem_bank[2772],db_odd.mem_bank[2773],db_even.mem_bank[2773],db_odd.mem_bank[2774],db_even.mem_bank[2774],db_odd.mem_bank[2775],db_even.mem_bank[2775],db_odd.mem_bank[2776],db_even.mem_bank[2776],db_odd.mem_bank[2777],db_even.mem_bank[2777],db_odd.mem_bank[2778],db_even.mem_bank[2778],db_odd.mem_bank[2779],db_even.mem_bank[2779],db_odd.mem_bank[2780],db_even.mem_bank[2780],db_odd.mem_bank[2781],db_even.mem_bank[2781],db_odd.mem_bank[2782],db_even.mem_bank[2782],db_odd.mem_bank[2783],db_even.mem_bank[2783],db_odd.mem_bank[2784],db_even.mem_bank[2784],db_odd.mem_bank[2785],db_even.mem_bank[2785],db_odd.mem_bank[2786],db_even.mem_bank[2786],db_odd.mem_bank[2787],db_even.mem_bank[2787],db_odd.mem_bank[2788],db_even.mem_bank[2788],db_odd.mem_bank[2789],db_even.mem_bank[2789],db_odd.mem_bank[2790],db_even.mem_bank[2790],db_odd.mem_bank[2791],db_even.mem_bank[2791],db_odd.mem_bank[2792],db_even.mem_bank[2792],db_odd.mem_bank[2793],db_even.mem_bank[2793],db_odd.mem_bank[2794],db_even.mem_bank[2794],db_odd.mem_bank[2795],db_even.mem_bank[2795],db_odd.mem_bank[2796],db_even.mem_bank[2796],db_odd.mem_bank[2797],db_even.mem_bank[2797],db_odd.mem_bank[2798],db_even.mem_bank[2798],db_odd.mem_bank[2799],db_even.mem_bank[2799],db_odd.mem_bank[2800],db_even.mem_bank[2800],db_odd.mem_bank[2801],db_even.mem_bank[2801],db_odd.mem_bank[2802],db_even.mem_bank[2802],db_odd.mem_bank[2803],db_even.mem_bank[2803],db_odd.mem_bank[2804],db_even.mem_bank[2804],db_odd.mem_bank[2805],db_even.mem_bank[2805],db_odd.mem_bank[2806],db_even.mem_bank[2806],db_odd.mem_bank[2807],db_even.mem_bank[2807],db_odd.mem_bank[2808],db_even.mem_bank[2808],db_odd.mem_bank[2809],db_even.mem_bank[2809],db_odd.mem_bank[2810],db_even.mem_bank[2810],db_odd.mem_bank[2811],db_even.mem_bank[2811],db_odd.mem_bank[2812],db_even.mem_bank[2812],db_odd.mem_bank[2813],db_even.mem_bank[2813],db_odd.mem_bank[2814],db_even.mem_bank[2814],db_odd.mem_bank[2815],db_even.mem_bank[2815],db_odd.mem_bank[2816],db_even.mem_bank[2816],db_odd.mem_bank[2817],db_even.mem_bank[2817],db_odd.mem_bank[2818],db_even.mem_bank[2818],db_odd.mem_bank[2819],db_even.mem_bank[2819],db_odd.mem_bank[2820],db_even.mem_bank[2820],db_odd.mem_bank[2821],db_even.mem_bank[2821],db_odd.mem_bank[2822],db_even.mem_bank[2822],db_odd.mem_bank[2823],db_even.mem_bank[2823],db_odd.mem_bank[2824],db_even.mem_bank[2824],db_odd.mem_bank[2825],db_even.mem_bank[2825],db_odd.mem_bank[2826],db_even.mem_bank[2826],db_odd.mem_bank[2827],db_even.mem_bank[2827],db_odd.mem_bank[2828],db_even.mem_bank[2828],db_odd.mem_bank[2829],db_even.mem_bank[2829],db_odd.mem_bank[2830],db_even.mem_bank[2830],db_odd.mem_bank[2831],db_even.mem_bank[2831],db_odd.mem_bank[2832],db_even.mem_bank[2832],db_odd.mem_bank[2833],db_even.mem_bank[2833],db_odd.mem_bank[2834],db_even.mem_bank[2834],db_odd.mem_bank[2835],db_even.mem_bank[2835],db_odd.mem_bank[2836],db_even.mem_bank[2836],db_odd.mem_bank[2837],db_even.mem_bank[2837],db_odd.mem_bank[2838],db_even.mem_bank[2838],db_odd.mem_bank[2839],db_even.mem_bank[2839],db_odd.mem_bank[2840],db_even.mem_bank[2840],db_odd.mem_bank[2841],db_even.mem_bank[2841],db_odd.mem_bank[2842],db_even.mem_bank[2842],db_odd.mem_bank[2843],db_even.mem_bank[2843],db_odd.mem_bank[2844],db_even.mem_bank[2844],db_odd.mem_bank[2845],db_even.mem_bank[2845],db_odd.mem_bank[2846],db_even.mem_bank[2846],db_odd.mem_bank[2847],db_even.mem_bank[2847],db_odd.mem_bank[2848],db_even.mem_bank[2848],db_odd.mem_bank[2849],db_even.mem_bank[2849],db_odd.mem_bank[2850],db_even.mem_bank[2850],db_odd.mem_bank[2851],db_even.mem_bank[2851],db_odd.mem_bank[2852],db_even.mem_bank[2852],db_odd.mem_bank[2853],db_even.mem_bank[2853],db_odd.mem_bank[2854],db_even.mem_bank[2854],db_odd.mem_bank[2855],db_even.mem_bank[2855],db_odd.mem_bank[2856],db_even.mem_bank[2856],db_odd.mem_bank[2857],db_even.mem_bank[2857],db_odd.mem_bank[2858],db_even.mem_bank[2858],db_odd.mem_bank[2859],db_even.mem_bank[2859],db_odd.mem_bank[2860],db_even.mem_bank[2860],db_odd.mem_bank[2861],db_even.mem_bank[2861],db_odd.mem_bank[2862],db_even.mem_bank[2862],db_odd.mem_bank[2863],db_even.mem_bank[2863],db_odd.mem_bank[2864],db_even.mem_bank[2864],db_odd.mem_bank[2865],db_even.mem_bank[2865],db_odd.mem_bank[2866],db_even.mem_bank[2866],db_odd.mem_bank[2867],db_even.mem_bank[2867],db_odd.mem_bank[2868],db_even.mem_bank[2868],db_odd.mem_bank[2869],db_even.mem_bank[2869],db_odd.mem_bank[2870],db_even.mem_bank[2870],db_odd.mem_bank[2871],db_even.mem_bank[2871],db_odd.mem_bank[2872],db_even.mem_bank[2872],db_odd.mem_bank[2873],db_even.mem_bank[2873],db_odd.mem_bank[2874],db_even.mem_bank[2874],db_odd.mem_bank[2875],db_even.mem_bank[2875],db_odd.mem_bank[2876],db_even.mem_bank[2876],db_odd.mem_bank[2877],db_even.mem_bank[2877],db_odd.mem_bank[2878],db_even.mem_bank[2878],db_odd.mem_bank[2879],db_even.mem_bank[2879],db_odd.mem_bank[2880],db_even.mem_bank[2880],db_odd.mem_bank[2881],db_even.mem_bank[2881],db_odd.mem_bank[2882],db_even.mem_bank[2882],db_odd.mem_bank[2883],db_even.mem_bank[2883],db_odd.mem_bank[2884],db_even.mem_bank[2884],db_odd.mem_bank[2885],db_even.mem_bank[2885],db_odd.mem_bank[2886],db_even.mem_bank[2886],db_odd.mem_bank[2887],db_even.mem_bank[2887],db_odd.mem_bank[2888],db_even.mem_bank[2888],db_odd.mem_bank[2889],db_even.mem_bank[2889],db_odd.mem_bank[2890],db_even.mem_bank[2890],db_odd.mem_bank[2891],db_even.mem_bank[2891],db_odd.mem_bank[2892],db_even.mem_bank[2892],db_odd.mem_bank[2893],db_even.mem_bank[2893],db_odd.mem_bank[2894],db_even.mem_bank[2894],db_odd.mem_bank[2895],db_even.mem_bank[2895],db_odd.mem_bank[2896],db_even.mem_bank[2896],db_odd.mem_bank[2897],db_even.mem_bank[2897],db_odd.mem_bank[2898],db_even.mem_bank[2898],db_odd.mem_bank[2899],db_even.mem_bank[2899],db_odd.mem_bank[2900],db_even.mem_bank[2900],db_odd.mem_bank[2901],db_even.mem_bank[2901],db_odd.mem_bank[2902],db_even.mem_bank[2902],db_odd.mem_bank[2903],db_even.mem_bank[2903],db_odd.mem_bank[2904],db_even.mem_bank[2904],db_odd.mem_bank[2905],db_even.mem_bank[2905],db_odd.mem_bank[2906],db_even.mem_bank[2906],db_odd.mem_bank[2907],db_even.mem_bank[2907],db_odd.mem_bank[2908],db_even.mem_bank[2908],db_odd.mem_bank[2909],db_even.mem_bank[2909],db_odd.mem_bank[2910],db_even.mem_bank[2910],db_odd.mem_bank[2911],db_even.mem_bank[2911],db_odd.mem_bank[2912],db_even.mem_bank[2912],db_odd.mem_bank[2913],db_even.mem_bank[2913],db_odd.mem_bank[2914],db_even.mem_bank[2914],db_odd.mem_bank[2915],db_even.mem_bank[2915],db_odd.mem_bank[2916],db_even.mem_bank[2916],db_odd.mem_bank[2917],db_even.mem_bank[2917],db_odd.mem_bank[2918],db_even.mem_bank[2918],db_odd.mem_bank[2919],db_even.mem_bank[2919],db_odd.mem_bank[2920],db_even.mem_bank[2920],db_odd.mem_bank[2921],db_even.mem_bank[2921],db_odd.mem_bank[2922],db_even.mem_bank[2922],db_odd.mem_bank[2923],db_even.mem_bank[2923],db_odd.mem_bank[2924],db_even.mem_bank[2924],db_odd.mem_bank[2925],db_even.mem_bank[2925],db_odd.mem_bank[2926],db_even.mem_bank[2926],db_odd.mem_bank[2927],db_even.mem_bank[2927],db_odd.mem_bank[2928],db_even.mem_bank[2928],db_odd.mem_bank[2929],db_even.mem_bank[2929],db_odd.mem_bank[2930],db_even.mem_bank[2930],db_odd.mem_bank[2931],db_even.mem_bank[2931],db_odd.mem_bank[2932],db_even.mem_bank[2932],db_odd.mem_bank[2933],db_even.mem_bank[2933],db_odd.mem_bank[2934],db_even.mem_bank[2934],db_odd.mem_bank[2935],db_even.mem_bank[2935],db_odd.mem_bank[2936],db_even.mem_bank[2936],db_odd.mem_bank[2937],db_even.mem_bank[2937],db_odd.mem_bank[2938],db_even.mem_bank[2938],db_odd.mem_bank[2939],db_even.mem_bank[2939],db_odd.mem_bank[2940],db_even.mem_bank[2940],db_odd.mem_bank[2941],db_even.mem_bank[2941],db_odd.mem_bank[2942],db_even.mem_bank[2942],db_odd.mem_bank[2943],db_even.mem_bank[2943],db_odd.mem_bank[2944],db_even.mem_bank[2944],db_odd.mem_bank[2945],db_even.mem_bank[2945],db_odd.mem_bank[2946],db_even.mem_bank[2946],db_odd.mem_bank[2947],db_even.mem_bank[2947],db_odd.mem_bank[2948],db_even.mem_bank[2948],db_odd.mem_bank[2949],db_even.mem_bank[2949],db_odd.mem_bank[2950],db_even.mem_bank[2950],db_odd.mem_bank[2951],db_even.mem_bank[2951],db_odd.mem_bank[2952],db_even.mem_bank[2952],db_odd.mem_bank[2953],db_even.mem_bank[2953],db_odd.mem_bank[2954],db_even.mem_bank[2954],db_odd.mem_bank[2955],db_even.mem_bank[2955],db_odd.mem_bank[2956],db_even.mem_bank[2956],db_odd.mem_bank[2957],db_even.mem_bank[2957],db_odd.mem_bank[2958],db_even.mem_bank[2958],db_odd.mem_bank[2959],db_even.mem_bank[2959],db_odd.mem_bank[2960],db_even.mem_bank[2960],db_odd.mem_bank[2961],db_even.mem_bank[2961],db_odd.mem_bank[2962],db_even.mem_bank[2962],db_odd.mem_bank[2963],db_even.mem_bank[2963],db_odd.mem_bank[2964],db_even.mem_bank[2964],db_odd.mem_bank[2965],db_even.mem_bank[2965],db_odd.mem_bank[2966],db_even.mem_bank[2966],db_odd.mem_bank[2967],db_even.mem_bank[2967],db_odd.mem_bank[2968],db_even.mem_bank[2968],db_odd.mem_bank[2969],db_even.mem_bank[2969],db_odd.mem_bank[2970],db_even.mem_bank[2970],db_odd.mem_bank[2971],db_even.mem_bank[2971],db_odd.mem_bank[2972],db_even.mem_bank[2972],db_odd.mem_bank[2973],db_even.mem_bank[2973],db_odd.mem_bank[2974],db_even.mem_bank[2974],db_odd.mem_bank[2975],db_even.mem_bank[2975],db_odd.mem_bank[2976],db_even.mem_bank[2976],db_odd.mem_bank[2977],db_even.mem_bank[2977],db_odd.mem_bank[2978],db_even.mem_bank[2978],db_odd.mem_bank[2979],db_even.mem_bank[2979],db_odd.mem_bank[2980],db_even.mem_bank[2980],db_odd.mem_bank[2981],db_even.mem_bank[2981],db_odd.mem_bank[2982],db_even.mem_bank[2982],db_odd.mem_bank[2983],db_even.mem_bank[2983],db_odd.mem_bank[2984],db_even.mem_bank[2984],db_odd.mem_bank[2985],db_even.mem_bank[2985],db_odd.mem_bank[2986],db_even.mem_bank[2986],db_odd.mem_bank[2987],db_even.mem_bank[2987],db_odd.mem_bank[2988],db_even.mem_bank[2988],db_odd.mem_bank[2989],db_even.mem_bank[2989],db_odd.mem_bank[2990],db_even.mem_bank[2990],db_odd.mem_bank[2991],db_even.mem_bank[2991],db_odd.mem_bank[2992],db_even.mem_bank[2992],db_odd.mem_bank[2993],db_even.mem_bank[2993],db_odd.mem_bank[2994],db_even.mem_bank[2994],db_odd.mem_bank[2995],db_even.mem_bank[2995],db_odd.mem_bank[2996],db_even.mem_bank[2996],db_odd.mem_bank[2997],db_even.mem_bank[2997],db_odd.mem_bank[2998],db_even.mem_bank[2998],db_odd.mem_bank[2999],db_even.mem_bank[2999],db_odd.mem_bank[3000],db_even.mem_bank[3000],db_odd.mem_bank[3001],db_even.mem_bank[3001],db_odd.mem_bank[3002],db_even.mem_bank[3002],db_odd.mem_bank[3003],db_even.mem_bank[3003],db_odd.mem_bank[3004],db_even.mem_bank[3004],db_odd.mem_bank[3005],db_even.mem_bank[3005],db_odd.mem_bank[3006],db_even.mem_bank[3006],db_odd.mem_bank[3007],db_even.mem_bank[3007],db_odd.mem_bank[3008],db_even.mem_bank[3008],db_odd.mem_bank[3009],db_even.mem_bank[3009],db_odd.mem_bank[3010],db_even.mem_bank[3010],db_odd.mem_bank[3011],db_even.mem_bank[3011],db_odd.mem_bank[3012],db_even.mem_bank[3012],db_odd.mem_bank[3013],db_even.mem_bank[3013],db_odd.mem_bank[3014],db_even.mem_bank[3014],db_odd.mem_bank[3015],db_even.mem_bank[3015],db_odd.mem_bank[3016],db_even.mem_bank[3016],db_odd.mem_bank[3017],db_even.mem_bank[3017],db_odd.mem_bank[3018],db_even.mem_bank[3018],db_odd.mem_bank[3019],db_even.mem_bank[3019],db_odd.mem_bank[3020],db_even.mem_bank[3020],db_odd.mem_bank[3021],db_even.mem_bank[3021],db_odd.mem_bank[3022],db_even.mem_bank[3022],db_odd.mem_bank[3023],db_even.mem_bank[3023],db_odd.mem_bank[3024],db_even.mem_bank[3024],db_odd.mem_bank[3025],db_even.mem_bank[3025],db_odd.mem_bank[3026],db_even.mem_bank[3026],db_odd.mem_bank[3027],db_even.mem_bank[3027],db_odd.mem_bank[3028],db_even.mem_bank[3028],db_odd.mem_bank[3029],db_even.mem_bank[3029],db_odd.mem_bank[3030],db_even.mem_bank[3030],db_odd.mem_bank[3031],db_even.mem_bank[3031],db_odd.mem_bank[3032],db_even.mem_bank[3032],db_odd.mem_bank[3033],db_even.mem_bank[3033],db_odd.mem_bank[3034],db_even.mem_bank[3034],db_odd.mem_bank[3035],db_even.mem_bank[3035],db_odd.mem_bank[3036],db_even.mem_bank[3036],db_odd.mem_bank[3037],db_even.mem_bank[3037],db_odd.mem_bank[3038],db_even.mem_bank[3038],db_odd.mem_bank[3039],db_even.mem_bank[3039],db_odd.mem_bank[3040],db_even.mem_bank[3040],db_odd.mem_bank[3041],db_even.mem_bank[3041],db_odd.mem_bank[3042],db_even.mem_bank[3042],db_odd.mem_bank[3043],db_even.mem_bank[3043],db_odd.mem_bank[3044],db_even.mem_bank[3044],db_odd.mem_bank[3045],db_even.mem_bank[3045],db_odd.mem_bank[3046],db_even.mem_bank[3046],db_odd.mem_bank[3047],db_even.mem_bank[3047],db_odd.mem_bank[3048],db_even.mem_bank[3048],db_odd.mem_bank[3049],db_even.mem_bank[3049],db_odd.mem_bank[3050],db_even.mem_bank[3050],db_odd.mem_bank[3051],db_even.mem_bank[3051],db_odd.mem_bank[3052],db_even.mem_bank[3052],db_odd.mem_bank[3053],db_even.mem_bank[3053],db_odd.mem_bank[3054],db_even.mem_bank[3054],db_odd.mem_bank[3055],db_even.mem_bank[3055],db_odd.mem_bank[3056],db_even.mem_bank[3056],db_odd.mem_bank[3057],db_even.mem_bank[3057],db_odd.mem_bank[3058],db_even.mem_bank[3058],db_odd.mem_bank[3059],db_even.mem_bank[3059],db_odd.mem_bank[3060],db_even.mem_bank[3060],db_odd.mem_bank[3061],db_even.mem_bank[3061],db_odd.mem_bank[3062],db_even.mem_bank[3062],db_odd.mem_bank[3063],db_even.mem_bank[3063],db_odd.mem_bank[3064],db_even.mem_bank[3064],db_odd.mem_bank[3065],db_even.mem_bank[3065],db_odd.mem_bank[3066],db_even.mem_bank[3066],db_odd.mem_bank[3067],db_even.mem_bank[3067],db_odd.mem_bank[3068],db_even.mem_bank[3068],db_odd.mem_bank[3069],db_even.mem_bank[3069],db_odd.mem_bank[3070],db_even.mem_bank[3070],db_odd.mem_bank[3071],db_even.mem_bank[3071],db_odd.mem_bank[3072],db_even.mem_bank[3072],db_odd.mem_bank[3073],db_even.mem_bank[3073],db_odd.mem_bank[3074],db_even.mem_bank[3074],db_odd.mem_bank[3075],db_even.mem_bank[3075],db_odd.mem_bank[3076],db_even.mem_bank[3076],db_odd.mem_bank[3077],db_even.mem_bank[3077],db_odd.mem_bank[3078],db_even.mem_bank[3078],db_odd.mem_bank[3079],db_even.mem_bank[3079],db_odd.mem_bank[3080],db_even.mem_bank[3080],db_odd.mem_bank[3081],db_even.mem_bank[3081],db_odd.mem_bank[3082],db_even.mem_bank[3082],db_odd.mem_bank[3083],db_even.mem_bank[3083],db_odd.mem_bank[3084],db_even.mem_bank[3084],db_odd.mem_bank[3085],db_even.mem_bank[3085],db_odd.mem_bank[3086],db_even.mem_bank[3086],db_odd.mem_bank[3087],db_even.mem_bank[3087],db_odd.mem_bank[3088],db_even.mem_bank[3088],db_odd.mem_bank[3089],db_even.mem_bank[3089],db_odd.mem_bank[3090],db_even.mem_bank[3090],db_odd.mem_bank[3091],db_even.mem_bank[3091],db_odd.mem_bank[3092],db_even.mem_bank[3092],db_odd.mem_bank[3093],db_even.mem_bank[3093],db_odd.mem_bank[3094],db_even.mem_bank[3094],db_odd.mem_bank[3095],db_even.mem_bank[3095],db_odd.mem_bank[3096],db_even.mem_bank[3096],db_odd.mem_bank[3097],db_even.mem_bank[3097],db_odd.mem_bank[3098],db_even.mem_bank[3098],db_odd.mem_bank[3099],db_even.mem_bank[3099],db_odd.mem_bank[3100],db_even.mem_bank[3100],db_odd.mem_bank[3101],db_even.mem_bank[3101],db_odd.mem_bank[3102],db_even.mem_bank[3102],db_odd.mem_bank[3103],db_even.mem_bank[3103],db_odd.mem_bank[3104],db_even.mem_bank[3104],db_odd.mem_bank[3105],db_even.mem_bank[3105],db_odd.mem_bank[3106],db_even.mem_bank[3106],db_odd.mem_bank[3107],db_even.mem_bank[3107],db_odd.mem_bank[3108],db_even.mem_bank[3108],db_odd.mem_bank[3109],db_even.mem_bank[3109],db_odd.mem_bank[3110],db_even.mem_bank[3110],db_odd.mem_bank[3111],db_even.mem_bank[3111],db_odd.mem_bank[3112],db_even.mem_bank[3112],db_odd.mem_bank[3113],db_even.mem_bank[3113],db_odd.mem_bank[3114],db_even.mem_bank[3114],db_odd.mem_bank[3115],db_even.mem_bank[3115],db_odd.mem_bank[3116],db_even.mem_bank[3116],db_odd.mem_bank[3117],db_even.mem_bank[3117],db_odd.mem_bank[3118],db_even.mem_bank[3118],db_odd.mem_bank[3119],db_even.mem_bank[3119],db_odd.mem_bank[3120],db_even.mem_bank[3120],db_odd.mem_bank[3121],db_even.mem_bank[3121],db_odd.mem_bank[3122],db_even.mem_bank[3122],db_odd.mem_bank[3123],db_even.mem_bank[3123],db_odd.mem_bank[3124],db_even.mem_bank[3124],db_odd.mem_bank[3125],db_even.mem_bank[3125],db_odd.mem_bank[3126],db_even.mem_bank[3126],db_odd.mem_bank[3127],db_even.mem_bank[3127],db_odd.mem_bank[3128],db_even.mem_bank[3128],db_odd.mem_bank[3129],db_even.mem_bank[3129],db_odd.mem_bank[3130],db_even.mem_bank[3130],db_odd.mem_bank[3131],db_even.mem_bank[3131],db_odd.mem_bank[3132],db_even.mem_bank[3132],db_odd.mem_bank[3133],db_even.mem_bank[3133],db_odd.mem_bank[3134],db_even.mem_bank[3134],db_odd.mem_bank[3135],db_even.mem_bank[3135],db_odd.mem_bank[3136],db_even.mem_bank[3136],db_odd.mem_bank[3137],db_even.mem_bank[3137],db_odd.mem_bank[3138],db_even.mem_bank[3138],db_odd.mem_bank[3139],db_even.mem_bank[3139],db_odd.mem_bank[3140],db_even.mem_bank[3140],db_odd.mem_bank[3141],db_even.mem_bank[3141],db_odd.mem_bank[3142],db_even.mem_bank[3142],db_odd.mem_bank[3143],db_even.mem_bank[3143],db_odd.mem_bank[3144],db_even.mem_bank[3144],db_odd.mem_bank[3145],db_even.mem_bank[3145],db_odd.mem_bank[3146],db_even.mem_bank[3146],db_odd.mem_bank[3147],db_even.mem_bank[3147],db_odd.mem_bank[3148],db_even.mem_bank[3148],db_odd.mem_bank[3149],db_even.mem_bank[3149],db_odd.mem_bank[3150],db_even.mem_bank[3150],db_odd.mem_bank[3151],db_even.mem_bank[3151],db_odd.mem_bank[3152],db_even.mem_bank[3152],db_odd.mem_bank[3153],db_even.mem_bank[3153],db_odd.mem_bank[3154],db_even.mem_bank[3154],db_odd.mem_bank[3155],db_even.mem_bank[3155],db_odd.mem_bank[3156],db_even.mem_bank[3156],db_odd.mem_bank[3157],db_even.mem_bank[3157],db_odd.mem_bank[3158],db_even.mem_bank[3158],db_odd.mem_bank[3159],db_even.mem_bank[3159],db_odd.mem_bank[3160],db_even.mem_bank[3160],db_odd.mem_bank[3161],db_even.mem_bank[3161],db_odd.mem_bank[3162],db_even.mem_bank[3162],db_odd.mem_bank[3163],db_even.mem_bank[3163],db_odd.mem_bank[3164],db_even.mem_bank[3164],db_odd.mem_bank[3165],db_even.mem_bank[3165],db_odd.mem_bank[3166],db_even.mem_bank[3166],db_odd.mem_bank[3167],db_even.mem_bank[3167],db_odd.mem_bank[3168],db_even.mem_bank[3168],db_odd.mem_bank[3169],db_even.mem_bank[3169],db_odd.mem_bank[3170],db_even.mem_bank[3170],db_odd.mem_bank[3171],db_even.mem_bank[3171],db_odd.mem_bank[3172],db_even.mem_bank[3172],db_odd.mem_bank[3173],db_even.mem_bank[3173],db_odd.mem_bank[3174],db_even.mem_bank[3174],db_odd.mem_bank[3175],db_even.mem_bank[3175],db_odd.mem_bank[3176],db_even.mem_bank[3176],db_odd.mem_bank[3177],db_even.mem_bank[3177],db_odd.mem_bank[3178],db_even.mem_bank[3178],db_odd.mem_bank[3179],db_even.mem_bank[3179],db_odd.mem_bank[3180],db_even.mem_bank[3180],db_odd.mem_bank[3181],db_even.mem_bank[3181],db_odd.mem_bank[3182],db_even.mem_bank[3182],db_odd.mem_bank[3183],db_even.mem_bank[3183],db_odd.mem_bank[3184],db_even.mem_bank[3184],db_odd.mem_bank[3185],db_even.mem_bank[3185],db_odd.mem_bank[3186],db_even.mem_bank[3186],db_odd.mem_bank[3187],db_even.mem_bank[3187],db_odd.mem_bank[3188],db_even.mem_bank[3188],db_odd.mem_bank[3189],db_even.mem_bank[3189],db_odd.mem_bank[3190],db_even.mem_bank[3190],db_odd.mem_bank[3191],db_even.mem_bank[3191],db_odd.mem_bank[3192],db_even.mem_bank[3192],db_odd.mem_bank[3193],db_even.mem_bank[3193],db_odd.mem_bank[3194],db_even.mem_bank[3194],db_odd.mem_bank[3195],db_even.mem_bank[3195],db_odd.mem_bank[3196],db_even.mem_bank[3196],db_odd.mem_bank[3197],db_even.mem_bank[3197],db_odd.mem_bank[3198],db_even.mem_bank[3198],db_odd.mem_bank[3199],db_even.mem_bank[3199],db_odd.mem_bank[3200],db_even.mem_bank[3200],db_odd.mem_bank[3201],db_even.mem_bank[3201],db_odd.mem_bank[3202],db_even.mem_bank[3202],db_odd.mem_bank[3203],db_even.mem_bank[3203],db_odd.mem_bank[3204],db_even.mem_bank[3204],db_odd.mem_bank[3205],db_even.mem_bank[3205],db_odd.mem_bank[3206],db_even.mem_bank[3206],db_odd.mem_bank[3207],db_even.mem_bank[3207],db_odd.mem_bank[3208],db_even.mem_bank[3208],db_odd.mem_bank[3209],db_even.mem_bank[3209],db_odd.mem_bank[3210],db_even.mem_bank[3210],db_odd.mem_bank[3211],db_even.mem_bank[3211],db_odd.mem_bank[3212],db_even.mem_bank[3212],db_odd.mem_bank[3213],db_even.mem_bank[3213],db_odd.mem_bank[3214],db_even.mem_bank[3214],db_odd.mem_bank[3215],db_even.mem_bank[3215],db_odd.mem_bank[3216],db_even.mem_bank[3216],db_odd.mem_bank[3217],db_even.mem_bank[3217],db_odd.mem_bank[3218],db_even.mem_bank[3218],db_odd.mem_bank[3219],db_even.mem_bank[3219],db_odd.mem_bank[3220],db_even.mem_bank[3220],db_odd.mem_bank[3221],db_even.mem_bank[3221],db_odd.mem_bank[3222],db_even.mem_bank[3222],db_odd.mem_bank[3223],db_even.mem_bank[3223],db_odd.mem_bank[3224],db_even.mem_bank[3224],db_odd.mem_bank[3225],db_even.mem_bank[3225],db_odd.mem_bank[3226],db_even.mem_bank[3226],db_odd.mem_bank[3227],db_even.mem_bank[3227],db_odd.mem_bank[3228],db_even.mem_bank[3228],db_odd.mem_bank[3229],db_even.mem_bank[3229],db_odd.mem_bank[3230],db_even.mem_bank[3230],db_odd.mem_bank[3231],db_even.mem_bank[3231],db_odd.mem_bank[3232],db_even.mem_bank[3232],db_odd.mem_bank[3233],db_even.mem_bank[3233],db_odd.mem_bank[3234],db_even.mem_bank[3234],db_odd.mem_bank[3235],db_even.mem_bank[3235],db_odd.mem_bank[3236],db_even.mem_bank[3236],db_odd.mem_bank[3237],db_even.mem_bank[3237],db_odd.mem_bank[3238],db_even.mem_bank[3238],db_odd.mem_bank[3239],db_even.mem_bank[3239],db_odd.mem_bank[3240],db_even.mem_bank[3240],db_odd.mem_bank[3241],db_even.mem_bank[3241],db_odd.mem_bank[3242],db_even.mem_bank[3242],db_odd.mem_bank[3243],db_even.mem_bank[3243],db_odd.mem_bank[3244],db_even.mem_bank[3244],db_odd.mem_bank[3245],db_even.mem_bank[3245],db_odd.mem_bank[3246],db_even.mem_bank[3246],db_odd.mem_bank[3247],db_even.mem_bank[3247],db_odd.mem_bank[3248],db_even.mem_bank[3248],db_odd.mem_bank[3249],db_even.mem_bank[3249],db_odd.mem_bank[3250],db_even.mem_bank[3250],db_odd.mem_bank[3251],db_even.mem_bank[3251],db_odd.mem_bank[3252],db_even.mem_bank[3252],db_odd.mem_bank[3253],db_even.mem_bank[3253],db_odd.mem_bank[3254],db_even.mem_bank[3254],db_odd.mem_bank[3255],db_even.mem_bank[3255],db_odd.mem_bank[3256],db_even.mem_bank[3256],db_odd.mem_bank[3257],db_even.mem_bank[3257],db_odd.mem_bank[3258],db_even.mem_bank[3258],db_odd.mem_bank[3259],db_even.mem_bank[3259],db_odd.mem_bank[3260],db_even.mem_bank[3260],db_odd.mem_bank[3261],db_even.mem_bank[3261],db_odd.mem_bank[3262],db_even.mem_bank[3262],db_odd.mem_bank[3263],db_even.mem_bank[3263],db_odd.mem_bank[3264],db_even.mem_bank[3264],db_odd.mem_bank[3265],db_even.mem_bank[3265],db_odd.mem_bank[3266],db_even.mem_bank[3266],db_odd.mem_bank[3267],db_even.mem_bank[3267],db_odd.mem_bank[3268],db_even.mem_bank[3268],db_odd.mem_bank[3269],db_even.mem_bank[3269],db_odd.mem_bank[3270],db_even.mem_bank[3270],db_odd.mem_bank[3271],db_even.mem_bank[3271],db_odd.mem_bank[3272],db_even.mem_bank[3272],db_odd.mem_bank[3273],db_even.mem_bank[3273],db_odd.mem_bank[3274],db_even.mem_bank[3274],db_odd.mem_bank[3275],db_even.mem_bank[3275],db_odd.mem_bank[3276],db_even.mem_bank[3276],db_odd.mem_bank[3277],db_even.mem_bank[3277],db_odd.mem_bank[3278],db_even.mem_bank[3278],db_odd.mem_bank[3279],db_even.mem_bank[3279],db_odd.mem_bank[3280],db_even.mem_bank[3280],db_odd.mem_bank[3281],db_even.mem_bank[3281],db_odd.mem_bank[3282],db_even.mem_bank[3282],db_odd.mem_bank[3283],db_even.mem_bank[3283],db_odd.mem_bank[3284],db_even.mem_bank[3284],db_odd.mem_bank[3285],db_even.mem_bank[3285],db_odd.mem_bank[3286],db_even.mem_bank[3286],db_odd.mem_bank[3287],db_even.mem_bank[3287],db_odd.mem_bank[3288],db_even.mem_bank[3288],db_odd.mem_bank[3289],db_even.mem_bank[3289],db_odd.mem_bank[3290],db_even.mem_bank[3290],db_odd.mem_bank[3291],db_even.mem_bank[3291],db_odd.mem_bank[3292],db_even.mem_bank[3292],db_odd.mem_bank[3293],db_even.mem_bank[3293],db_odd.mem_bank[3294],db_even.mem_bank[3294],db_odd.mem_bank[3295],db_even.mem_bank[3295],db_odd.mem_bank[3296],db_even.mem_bank[3296],db_odd.mem_bank[3297],db_even.mem_bank[3297],db_odd.mem_bank[3298],db_even.mem_bank[3298],db_odd.mem_bank[3299],db_even.mem_bank[3299],db_odd.mem_bank[3300],db_even.mem_bank[3300],db_odd.mem_bank[3301],db_even.mem_bank[3301],db_odd.mem_bank[3302],db_even.mem_bank[3302],db_odd.mem_bank[3303],db_even.mem_bank[3303],db_odd.mem_bank[3304],db_even.mem_bank[3304],db_odd.mem_bank[3305],db_even.mem_bank[3305],db_odd.mem_bank[3306],db_even.mem_bank[3306],db_odd.mem_bank[3307],db_even.mem_bank[3307],db_odd.mem_bank[3308],db_even.mem_bank[3308],db_odd.mem_bank[3309],db_even.mem_bank[3309],db_odd.mem_bank[3310],db_even.mem_bank[3310],db_odd.mem_bank[3311],db_even.mem_bank[3311],db_odd.mem_bank[3312],db_even.mem_bank[3312],db_odd.mem_bank[3313],db_even.mem_bank[3313],db_odd.mem_bank[3314],db_even.mem_bank[3314],db_odd.mem_bank[3315],db_even.mem_bank[3315],db_odd.mem_bank[3316],db_even.mem_bank[3316],db_odd.mem_bank[3317],db_even.mem_bank[3317],db_odd.mem_bank[3318],db_even.mem_bank[3318],db_odd.mem_bank[3319],db_even.mem_bank[3319],db_odd.mem_bank[3320],db_even.mem_bank[3320],db_odd.mem_bank[3321],db_even.mem_bank[3321],db_odd.mem_bank[3322],db_even.mem_bank[3322],db_odd.mem_bank[3323],db_even.mem_bank[3323],db_odd.mem_bank[3324],db_even.mem_bank[3324],db_odd.mem_bank[3325],db_even.mem_bank[3325],db_odd.mem_bank[3326],db_even.mem_bank[3326],db_odd.mem_bank[3327],db_even.mem_bank[3327],db_odd.mem_bank[3328],db_even.mem_bank[3328],db_odd.mem_bank[3329],db_even.mem_bank[3329],db_odd.mem_bank[3330],db_even.mem_bank[3330],db_odd.mem_bank[3331],db_even.mem_bank[3331],db_odd.mem_bank[3332],db_even.mem_bank[3332],db_odd.mem_bank[3333],db_even.mem_bank[3333],db_odd.mem_bank[3334],db_even.mem_bank[3334],db_odd.mem_bank[3335],db_even.mem_bank[3335],db_odd.mem_bank[3336],db_even.mem_bank[3336],db_odd.mem_bank[3337],db_even.mem_bank[3337],db_odd.mem_bank[3338],db_even.mem_bank[3338],db_odd.mem_bank[3339],db_even.mem_bank[3339],db_odd.mem_bank[3340],db_even.mem_bank[3340],db_odd.mem_bank[3341],db_even.mem_bank[3341],db_odd.mem_bank[3342],db_even.mem_bank[3342],db_odd.mem_bank[3343],db_even.mem_bank[3343],db_odd.mem_bank[3344],db_even.mem_bank[3344],db_odd.mem_bank[3345],db_even.mem_bank[3345],db_odd.mem_bank[3346],db_even.mem_bank[3346],db_odd.mem_bank[3347],db_even.mem_bank[3347],db_odd.mem_bank[3348],db_even.mem_bank[3348],db_odd.mem_bank[3349],db_even.mem_bank[3349],db_odd.mem_bank[3350],db_even.mem_bank[3350],db_odd.mem_bank[3351],db_even.mem_bank[3351],db_odd.mem_bank[3352],db_even.mem_bank[3352],db_odd.mem_bank[3353],db_even.mem_bank[3353],db_odd.mem_bank[3354],db_even.mem_bank[3354],db_odd.mem_bank[3355],db_even.mem_bank[3355],db_odd.mem_bank[3356],db_even.mem_bank[3356],db_odd.mem_bank[3357],db_even.mem_bank[3357],db_odd.mem_bank[3358],db_even.mem_bank[3358],db_odd.mem_bank[3359],db_even.mem_bank[3359],db_odd.mem_bank[3360],db_even.mem_bank[3360],db_odd.mem_bank[3361],db_even.mem_bank[3361],db_odd.mem_bank[3362],db_even.mem_bank[3362],db_odd.mem_bank[3363],db_even.mem_bank[3363],db_odd.mem_bank[3364],db_even.mem_bank[3364],db_odd.mem_bank[3365],db_even.mem_bank[3365],db_odd.mem_bank[3366],db_even.mem_bank[3366],db_odd.mem_bank[3367],db_even.mem_bank[3367],db_odd.mem_bank[3368],db_even.mem_bank[3368],db_odd.mem_bank[3369],db_even.mem_bank[3369],db_odd.mem_bank[3370],db_even.mem_bank[3370],db_odd.mem_bank[3371],db_even.mem_bank[3371],db_odd.mem_bank[3372],db_even.mem_bank[3372],db_odd.mem_bank[3373],db_even.mem_bank[3373],db_odd.mem_bank[3374],db_even.mem_bank[3374],db_odd.mem_bank[3375],db_even.mem_bank[3375],db_odd.mem_bank[3376],db_even.mem_bank[3376],db_odd.mem_bank[3377],db_even.mem_bank[3377],db_odd.mem_bank[3378],db_even.mem_bank[3378],db_odd.mem_bank[3379],db_even.mem_bank[3379],db_odd.mem_bank[3380],db_even.mem_bank[3380],db_odd.mem_bank[3381],db_even.mem_bank[3381],db_odd.mem_bank[3382],db_even.mem_bank[3382],db_odd.mem_bank[3383],db_even.mem_bank[3383],db_odd.mem_bank[3384],db_even.mem_bank[3384],db_odd.mem_bank[3385],db_even.mem_bank[3385],db_odd.mem_bank[3386],db_even.mem_bank[3386],db_odd.mem_bank[3387],db_even.mem_bank[3387],db_odd.mem_bank[3388],db_even.mem_bank[3388],db_odd.mem_bank[3389],db_even.mem_bank[3389],db_odd.mem_bank[3390],db_even.mem_bank[3390],db_odd.mem_bank[3391],db_even.mem_bank[3391],db_odd.mem_bank[3392],db_even.mem_bank[3392],db_odd.mem_bank[3393],db_even.mem_bank[3393],db_odd.mem_bank[3394],db_even.mem_bank[3394],db_odd.mem_bank[3395],db_even.mem_bank[3395],db_odd.mem_bank[3396],db_even.mem_bank[3396],db_odd.mem_bank[3397],db_even.mem_bank[3397],db_odd.mem_bank[3398],db_even.mem_bank[3398],db_odd.mem_bank[3399],db_even.mem_bank[3399],db_odd.mem_bank[3400],db_even.mem_bank[3400],db_odd.mem_bank[3401],db_even.mem_bank[3401],db_odd.mem_bank[3402],db_even.mem_bank[3402],db_odd.mem_bank[3403],db_even.mem_bank[3403],db_odd.mem_bank[3404],db_even.mem_bank[3404],db_odd.mem_bank[3405],db_even.mem_bank[3405],db_odd.mem_bank[3406],db_even.mem_bank[3406],db_odd.mem_bank[3407],db_even.mem_bank[3407],db_odd.mem_bank[3408],db_even.mem_bank[3408],db_odd.mem_bank[3409],db_even.mem_bank[3409],db_odd.mem_bank[3410],db_even.mem_bank[3410],db_odd.mem_bank[3411],db_even.mem_bank[3411],db_odd.mem_bank[3412],db_even.mem_bank[3412],db_odd.mem_bank[3413],db_even.mem_bank[3413],db_odd.mem_bank[3414],db_even.mem_bank[3414],db_odd.mem_bank[3415],db_even.mem_bank[3415],db_odd.mem_bank[3416],db_even.mem_bank[3416],db_odd.mem_bank[3417],db_even.mem_bank[3417],db_odd.mem_bank[3418],db_even.mem_bank[3418],db_odd.mem_bank[3419],db_even.mem_bank[3419],db_odd.mem_bank[3420],db_even.mem_bank[3420],db_odd.mem_bank[3421],db_even.mem_bank[3421],db_odd.mem_bank[3422],db_even.mem_bank[3422],db_odd.mem_bank[3423],db_even.mem_bank[3423],db_odd.mem_bank[3424],db_even.mem_bank[3424],db_odd.mem_bank[3425],db_even.mem_bank[3425],db_odd.mem_bank[3426],db_even.mem_bank[3426],db_odd.mem_bank[3427],db_even.mem_bank[3427],db_odd.mem_bank[3428],db_even.mem_bank[3428],db_odd.mem_bank[3429],db_even.mem_bank[3429],db_odd.mem_bank[3430],db_even.mem_bank[3430],db_odd.mem_bank[3431],db_even.mem_bank[3431],db_odd.mem_bank[3432],db_even.mem_bank[3432],db_odd.mem_bank[3433],db_even.mem_bank[3433],db_odd.mem_bank[3434],db_even.mem_bank[3434],db_odd.mem_bank[3435],db_even.mem_bank[3435],db_odd.mem_bank[3436],db_even.mem_bank[3436],db_odd.mem_bank[3437],db_even.mem_bank[3437],db_odd.mem_bank[3438],db_even.mem_bank[3438],db_odd.mem_bank[3439],db_even.mem_bank[3439],db_odd.mem_bank[3440],db_even.mem_bank[3440],db_odd.mem_bank[3441],db_even.mem_bank[3441],db_odd.mem_bank[3442],db_even.mem_bank[3442],db_odd.mem_bank[3443],db_even.mem_bank[3443],db_odd.mem_bank[3444],db_even.mem_bank[3444],db_odd.mem_bank[3445],db_even.mem_bank[3445],db_odd.mem_bank[3446],db_even.mem_bank[3446],db_odd.mem_bank[3447],db_even.mem_bank[3447],db_odd.mem_bank[3448],db_even.mem_bank[3448],db_odd.mem_bank[3449],db_even.mem_bank[3449],db_odd.mem_bank[3450],db_even.mem_bank[3450],db_odd.mem_bank[3451],db_even.mem_bank[3451],db_odd.mem_bank[3452],db_even.mem_bank[3452],db_odd.mem_bank[3453],db_even.mem_bank[3453],db_odd.mem_bank[3454],db_even.mem_bank[3454],db_odd.mem_bank[3455],db_even.mem_bank[3455],db_odd.mem_bank[3456],db_even.mem_bank[3456],db_odd.mem_bank[3457],db_even.mem_bank[3457],db_odd.mem_bank[3458],db_even.mem_bank[3458],db_odd.mem_bank[3459],db_even.mem_bank[3459],db_odd.mem_bank[3460],db_even.mem_bank[3460],db_odd.mem_bank[3461],db_even.mem_bank[3461],db_odd.mem_bank[3462],db_even.mem_bank[3462],db_odd.mem_bank[3463],db_even.mem_bank[3463],db_odd.mem_bank[3464],db_even.mem_bank[3464],db_odd.mem_bank[3465],db_even.mem_bank[3465],db_odd.mem_bank[3466],db_even.mem_bank[3466],db_odd.mem_bank[3467],db_even.mem_bank[3467],db_odd.mem_bank[3468],db_even.mem_bank[3468],db_odd.mem_bank[3469],db_even.mem_bank[3469],db_odd.mem_bank[3470],db_even.mem_bank[3470],db_odd.mem_bank[3471],db_even.mem_bank[3471],db_odd.mem_bank[3472],db_even.mem_bank[3472],db_odd.mem_bank[3473],db_even.mem_bank[3473],db_odd.mem_bank[3474],db_even.mem_bank[3474],db_odd.mem_bank[3475],db_even.mem_bank[3475],db_odd.mem_bank[3476],db_even.mem_bank[3476],db_odd.mem_bank[3477],db_even.mem_bank[3477],db_odd.mem_bank[3478],db_even.mem_bank[3478],db_odd.mem_bank[3479],db_even.mem_bank[3479],db_odd.mem_bank[3480],db_even.mem_bank[3480],db_odd.mem_bank[3481],db_even.mem_bank[3481],db_odd.mem_bank[3482],db_even.mem_bank[3482],db_odd.mem_bank[3483],db_even.mem_bank[3483],db_odd.mem_bank[3484],db_even.mem_bank[3484],db_odd.mem_bank[3485],db_even.mem_bank[3485],db_odd.mem_bank[3486],db_even.mem_bank[3486],db_odd.mem_bank[3487],db_even.mem_bank[3487],db_odd.mem_bank[3488],db_even.mem_bank[3488],db_odd.mem_bank[3489],db_even.mem_bank[3489],db_odd.mem_bank[3490],db_even.mem_bank[3490],db_odd.mem_bank[3491],db_even.mem_bank[3491],db_odd.mem_bank[3492],db_even.mem_bank[3492],db_odd.mem_bank[3493],db_even.mem_bank[3493],db_odd.mem_bank[3494],db_even.mem_bank[3494],db_odd.mem_bank[3495],db_even.mem_bank[3495],db_odd.mem_bank[3496],db_even.mem_bank[3496],db_odd.mem_bank[3497],db_even.mem_bank[3497],db_odd.mem_bank[3498],db_even.mem_bank[3498],db_odd.mem_bank[3499],db_even.mem_bank[3499],db_odd.mem_bank[3500],db_even.mem_bank[3500],db_odd.mem_bank[3501],db_even.mem_bank[3501],db_odd.mem_bank[3502],db_even.mem_bank[3502],db_odd.mem_bank[3503],db_even.mem_bank[3503],db_odd.mem_bank[3504],db_even.mem_bank[3504],db_odd.mem_bank[3505],db_even.mem_bank[3505],db_odd.mem_bank[3506],db_even.mem_bank[3506],db_odd.mem_bank[3507],db_even.mem_bank[3507],db_odd.mem_bank[3508],db_even.mem_bank[3508],db_odd.mem_bank[3509],db_even.mem_bank[3509],db_odd.mem_bank[3510],db_even.mem_bank[3510],db_odd.mem_bank[3511],db_even.mem_bank[3511],db_odd.mem_bank[3512],db_even.mem_bank[3512],db_odd.mem_bank[3513],db_even.mem_bank[3513],db_odd.mem_bank[3514],db_even.mem_bank[3514],db_odd.mem_bank[3515],db_even.mem_bank[3515],db_odd.mem_bank[3516],db_even.mem_bank[3516],db_odd.mem_bank[3517],db_even.mem_bank[3517],db_odd.mem_bank[3518],db_even.mem_bank[3518],db_odd.mem_bank[3519],db_even.mem_bank[3519],db_odd.mem_bank[3520],db_even.mem_bank[3520],db_odd.mem_bank[3521],db_even.mem_bank[3521],db_odd.mem_bank[3522],db_even.mem_bank[3522],db_odd.mem_bank[3523],db_even.mem_bank[3523],db_odd.mem_bank[3524],db_even.mem_bank[3524],db_odd.mem_bank[3525],db_even.mem_bank[3525],db_odd.mem_bank[3526],db_even.mem_bank[3526],db_odd.mem_bank[3527],db_even.mem_bank[3527],db_odd.mem_bank[3528],db_even.mem_bank[3528],db_odd.mem_bank[3529],db_even.mem_bank[3529],db_odd.mem_bank[3530],db_even.mem_bank[3530],db_odd.mem_bank[3531],db_even.mem_bank[3531],db_odd.mem_bank[3532],db_even.mem_bank[3532],db_odd.mem_bank[3533],db_even.mem_bank[3533],db_odd.mem_bank[3534],db_even.mem_bank[3534],db_odd.mem_bank[3535],db_even.mem_bank[3535],db_odd.mem_bank[3536],db_even.mem_bank[3536],db_odd.mem_bank[3537],db_even.mem_bank[3537],db_odd.mem_bank[3538],db_even.mem_bank[3538],db_odd.mem_bank[3539],db_even.mem_bank[3539],db_odd.mem_bank[3540],db_even.mem_bank[3540],db_odd.mem_bank[3541],db_even.mem_bank[3541],db_odd.mem_bank[3542],db_even.mem_bank[3542],db_odd.mem_bank[3543],db_even.mem_bank[3543],db_odd.mem_bank[3544],db_even.mem_bank[3544],db_odd.mem_bank[3545],db_even.mem_bank[3545],db_odd.mem_bank[3546],db_even.mem_bank[3546],db_odd.mem_bank[3547],db_even.mem_bank[3547],db_odd.mem_bank[3548],db_even.mem_bank[3548],db_odd.mem_bank[3549],db_even.mem_bank[3549],db_odd.mem_bank[3550],db_even.mem_bank[3550],db_odd.mem_bank[3551],db_even.mem_bank[3551],db_odd.mem_bank[3552],db_even.mem_bank[3552],db_odd.mem_bank[3553],db_even.mem_bank[3553],db_odd.mem_bank[3554],db_even.mem_bank[3554],db_odd.mem_bank[3555],db_even.mem_bank[3555],db_odd.mem_bank[3556],db_even.mem_bank[3556],db_odd.mem_bank[3557],db_even.mem_bank[3557],db_odd.mem_bank[3558],db_even.mem_bank[3558],db_odd.mem_bank[3559],db_even.mem_bank[3559],db_odd.mem_bank[3560],db_even.mem_bank[3560],db_odd.mem_bank[3561],db_even.mem_bank[3561],db_odd.mem_bank[3562],db_even.mem_bank[3562],db_odd.mem_bank[3563],db_even.mem_bank[3563],db_odd.mem_bank[3564],db_even.mem_bank[3564],db_odd.mem_bank[3565],db_even.mem_bank[3565],db_odd.mem_bank[3566],db_even.mem_bank[3566],db_odd.mem_bank[3567],db_even.mem_bank[3567],db_odd.mem_bank[3568],db_even.mem_bank[3568],db_odd.mem_bank[3569],db_even.mem_bank[3569],db_odd.mem_bank[3570],db_even.mem_bank[3570],db_odd.mem_bank[3571],db_even.mem_bank[3571],db_odd.mem_bank[3572],db_even.mem_bank[3572],db_odd.mem_bank[3573],db_even.mem_bank[3573],db_odd.mem_bank[3574],db_even.mem_bank[3574],db_odd.mem_bank[3575],db_even.mem_bank[3575],db_odd.mem_bank[3576],db_even.mem_bank[3576],db_odd.mem_bank[3577],db_even.mem_bank[3577],db_odd.mem_bank[3578],db_even.mem_bank[3578],db_odd.mem_bank[3579],db_even.mem_bank[3579],db_odd.mem_bank[3580],db_even.mem_bank[3580],db_odd.mem_bank[3581],db_even.mem_bank[3581],db_odd.mem_bank[3582],db_even.mem_bank[3582],db_odd.mem_bank[3583],db_even.mem_bank[3583],db_odd.mem_bank[3584],db_even.mem_bank[3584],db_odd.mem_bank[3585],db_even.mem_bank[3585],db_odd.mem_bank[3586],db_even.mem_bank[3586],db_odd.mem_bank[3587],db_even.mem_bank[3587],db_odd.mem_bank[3588],db_even.mem_bank[3588],db_odd.mem_bank[3589],db_even.mem_bank[3589],db_odd.mem_bank[3590],db_even.mem_bank[3590],db_odd.mem_bank[3591],db_even.mem_bank[3591],db_odd.mem_bank[3592],db_even.mem_bank[3592],db_odd.mem_bank[3593],db_even.mem_bank[3593],db_odd.mem_bank[3594],db_even.mem_bank[3594],db_odd.mem_bank[3595],db_even.mem_bank[3595],db_odd.mem_bank[3596],db_even.mem_bank[3596],db_odd.mem_bank[3597],db_even.mem_bank[3597],db_odd.mem_bank[3598],db_even.mem_bank[3598],db_odd.mem_bank[3599],db_even.mem_bank[3599],db_odd.mem_bank[3600],db_even.mem_bank[3600],db_odd.mem_bank[3601],db_even.mem_bank[3601],db_odd.mem_bank[3602],db_even.mem_bank[3602],db_odd.mem_bank[3603],db_even.mem_bank[3603],db_odd.mem_bank[3604],db_even.mem_bank[3604],db_odd.mem_bank[3605],db_even.mem_bank[3605],db_odd.mem_bank[3606],db_even.mem_bank[3606],db_odd.mem_bank[3607],db_even.mem_bank[3607],db_odd.mem_bank[3608],db_even.mem_bank[3608],db_odd.mem_bank[3609],db_even.mem_bank[3609],db_odd.mem_bank[3610],db_even.mem_bank[3610],db_odd.mem_bank[3611],db_even.mem_bank[3611],db_odd.mem_bank[3612],db_even.mem_bank[3612],db_odd.mem_bank[3613],db_even.mem_bank[3613],db_odd.mem_bank[3614],db_even.mem_bank[3614],db_odd.mem_bank[3615],db_even.mem_bank[3615],db_odd.mem_bank[3616],db_even.mem_bank[3616],db_odd.mem_bank[3617],db_even.mem_bank[3617],db_odd.mem_bank[3618],db_even.mem_bank[3618],db_odd.mem_bank[3619],db_even.mem_bank[3619],db_odd.mem_bank[3620],db_even.mem_bank[3620],db_odd.mem_bank[3621],db_even.mem_bank[3621],db_odd.mem_bank[3622],db_even.mem_bank[3622],db_odd.mem_bank[3623],db_even.mem_bank[3623],db_odd.mem_bank[3624],db_even.mem_bank[3624],db_odd.mem_bank[3625],db_even.mem_bank[3625],db_odd.mem_bank[3626],db_even.mem_bank[3626],db_odd.mem_bank[3627],db_even.mem_bank[3627],db_odd.mem_bank[3628],db_even.mem_bank[3628],db_odd.mem_bank[3629],db_even.mem_bank[3629],db_odd.mem_bank[3630],db_even.mem_bank[3630],db_odd.mem_bank[3631],db_even.mem_bank[3631],db_odd.mem_bank[3632],db_even.mem_bank[3632],db_odd.mem_bank[3633],db_even.mem_bank[3633],db_odd.mem_bank[3634],db_even.mem_bank[3634],db_odd.mem_bank[3635],db_even.mem_bank[3635],db_odd.mem_bank[3636],db_even.mem_bank[3636],db_odd.mem_bank[3637],db_even.mem_bank[3637],db_odd.mem_bank[3638],db_even.mem_bank[3638],db_odd.mem_bank[3639],db_even.mem_bank[3639],db_odd.mem_bank[3640],db_even.mem_bank[3640],db_odd.mem_bank[3641],db_even.mem_bank[3641],db_odd.mem_bank[3642],db_even.mem_bank[3642],db_odd.mem_bank[3643],db_even.mem_bank[3643],db_odd.mem_bank[3644],db_even.mem_bank[3644],db_odd.mem_bank[3645],db_even.mem_bank[3645],db_odd.mem_bank[3646],db_even.mem_bank[3646],db_odd.mem_bank[3647],db_even.mem_bank[3647],db_odd.mem_bank[3648],db_even.mem_bank[3648],db_odd.mem_bank[3649],db_even.mem_bank[3649],db_odd.mem_bank[3650],db_even.mem_bank[3650],db_odd.mem_bank[3651],db_even.mem_bank[3651],db_odd.mem_bank[3652],db_even.mem_bank[3652],db_odd.mem_bank[3653],db_even.mem_bank[3653],db_odd.mem_bank[3654],db_even.mem_bank[3654],db_odd.mem_bank[3655],db_even.mem_bank[3655],db_odd.mem_bank[3656],db_even.mem_bank[3656],db_odd.mem_bank[3657],db_even.mem_bank[3657],db_odd.mem_bank[3658],db_even.mem_bank[3658],db_odd.mem_bank[3659],db_even.mem_bank[3659],db_odd.mem_bank[3660],db_even.mem_bank[3660],db_odd.mem_bank[3661],db_even.mem_bank[3661],db_odd.mem_bank[3662],db_even.mem_bank[3662],db_odd.mem_bank[3663],db_even.mem_bank[3663],db_odd.mem_bank[3664],db_even.mem_bank[3664],db_odd.mem_bank[3665],db_even.mem_bank[3665],db_odd.mem_bank[3666],db_even.mem_bank[3666],db_odd.mem_bank[3667],db_even.mem_bank[3667],db_odd.mem_bank[3668],db_even.mem_bank[3668],db_odd.mem_bank[3669],db_even.mem_bank[3669],db_odd.mem_bank[3670],db_even.mem_bank[3670],db_odd.mem_bank[3671],db_even.mem_bank[3671],db_odd.mem_bank[3672],db_even.mem_bank[3672],db_odd.mem_bank[3673],db_even.mem_bank[3673],db_odd.mem_bank[3674],db_even.mem_bank[3674],db_odd.mem_bank[3675],db_even.mem_bank[3675],db_odd.mem_bank[3676],db_even.mem_bank[3676],db_odd.mem_bank[3677],db_even.mem_bank[3677],db_odd.mem_bank[3678],db_even.mem_bank[3678],db_odd.mem_bank[3679],db_even.mem_bank[3679],db_odd.mem_bank[3680],db_even.mem_bank[3680],db_odd.mem_bank[3681],db_even.mem_bank[3681],db_odd.mem_bank[3682],db_even.mem_bank[3682],db_odd.mem_bank[3683],db_even.mem_bank[3683],db_odd.mem_bank[3684],db_even.mem_bank[3684],db_odd.mem_bank[3685],db_even.mem_bank[3685],db_odd.mem_bank[3686],db_even.mem_bank[3686],db_odd.mem_bank[3687],db_even.mem_bank[3687],db_odd.mem_bank[3688],db_even.mem_bank[3688],db_odd.mem_bank[3689],db_even.mem_bank[3689],db_odd.mem_bank[3690],db_even.mem_bank[3690],db_odd.mem_bank[3691],db_even.mem_bank[3691],db_odd.mem_bank[3692],db_even.mem_bank[3692],db_odd.mem_bank[3693],db_even.mem_bank[3693],db_odd.mem_bank[3694],db_even.mem_bank[3694],db_odd.mem_bank[3695],db_even.mem_bank[3695],db_odd.mem_bank[3696],db_even.mem_bank[3696],db_odd.mem_bank[3697],db_even.mem_bank[3697],db_odd.mem_bank[3698],db_even.mem_bank[3698],db_odd.mem_bank[3699],db_even.mem_bank[3699],db_odd.mem_bank[3700],db_even.mem_bank[3700],db_odd.mem_bank[3701],db_even.mem_bank[3701],db_odd.mem_bank[3702],db_even.mem_bank[3702],db_odd.mem_bank[3703],db_even.mem_bank[3703],db_odd.mem_bank[3704],db_even.mem_bank[3704],db_odd.mem_bank[3705],db_even.mem_bank[3705],db_odd.mem_bank[3706],db_even.mem_bank[3706],db_odd.mem_bank[3707],db_even.mem_bank[3707],db_odd.mem_bank[3708],db_even.mem_bank[3708],db_odd.mem_bank[3709],db_even.mem_bank[3709],db_odd.mem_bank[3710],db_even.mem_bank[3710],db_odd.mem_bank[3711],db_even.mem_bank[3711],db_odd.mem_bank[3712],db_even.mem_bank[3712],db_odd.mem_bank[3713],db_even.mem_bank[3713],db_odd.mem_bank[3714],db_even.mem_bank[3714],db_odd.mem_bank[3715],db_even.mem_bank[3715],db_odd.mem_bank[3716],db_even.mem_bank[3716],db_odd.mem_bank[3717],db_even.mem_bank[3717],db_odd.mem_bank[3718],db_even.mem_bank[3718],db_odd.mem_bank[3719],db_even.mem_bank[3719],db_odd.mem_bank[3720],db_even.mem_bank[3720],db_odd.mem_bank[3721],db_even.mem_bank[3721],db_odd.mem_bank[3722],db_even.mem_bank[3722],db_odd.mem_bank[3723],db_even.mem_bank[3723],db_odd.mem_bank[3724],db_even.mem_bank[3724],db_odd.mem_bank[3725],db_even.mem_bank[3725],db_odd.mem_bank[3726],db_even.mem_bank[3726],db_odd.mem_bank[3727],db_even.mem_bank[3727],db_odd.mem_bank[3728],db_even.mem_bank[3728],db_odd.mem_bank[3729],db_even.mem_bank[3729],db_odd.mem_bank[3730],db_even.mem_bank[3730],db_odd.mem_bank[3731],db_even.mem_bank[3731],db_odd.mem_bank[3732],db_even.mem_bank[3732],db_odd.mem_bank[3733],db_even.mem_bank[3733],db_odd.mem_bank[3734],db_even.mem_bank[3734],db_odd.mem_bank[3735],db_even.mem_bank[3735],db_odd.mem_bank[3736],db_even.mem_bank[3736],db_odd.mem_bank[3737],db_even.mem_bank[3737],db_odd.mem_bank[3738],db_even.mem_bank[3738],db_odd.mem_bank[3739],db_even.mem_bank[3739],db_odd.mem_bank[3740],db_even.mem_bank[3740],db_odd.mem_bank[3741],db_even.mem_bank[3741],db_odd.mem_bank[3742],db_even.mem_bank[3742],db_odd.mem_bank[3743],db_even.mem_bank[3743],db_odd.mem_bank[3744],db_even.mem_bank[3744],db_odd.mem_bank[3745],db_even.mem_bank[3745],db_odd.mem_bank[3746],db_even.mem_bank[3746],db_odd.mem_bank[3747],db_even.mem_bank[3747],db_odd.mem_bank[3748],db_even.mem_bank[3748],db_odd.mem_bank[3749],db_even.mem_bank[3749],db_odd.mem_bank[3750],db_even.mem_bank[3750],db_odd.mem_bank[3751],db_even.mem_bank[3751],db_odd.mem_bank[3752],db_even.mem_bank[3752],db_odd.mem_bank[3753],db_even.mem_bank[3753],db_odd.mem_bank[3754],db_even.mem_bank[3754],db_odd.mem_bank[3755],db_even.mem_bank[3755],db_odd.mem_bank[3756],db_even.mem_bank[3756],db_odd.mem_bank[3757],db_even.mem_bank[3757],db_odd.mem_bank[3758],db_even.mem_bank[3758],db_odd.mem_bank[3759],db_even.mem_bank[3759],db_odd.mem_bank[3760],db_even.mem_bank[3760],db_odd.mem_bank[3761],db_even.mem_bank[3761],db_odd.mem_bank[3762],db_even.mem_bank[3762],db_odd.mem_bank[3763],db_even.mem_bank[3763],db_odd.mem_bank[3764],db_even.mem_bank[3764],db_odd.mem_bank[3765],db_even.mem_bank[3765],db_odd.mem_bank[3766],db_even.mem_bank[3766],db_odd.mem_bank[3767],db_even.mem_bank[3767],db_odd.mem_bank[3768],db_even.mem_bank[3768],db_odd.mem_bank[3769],db_even.mem_bank[3769],db_odd.mem_bank[3770],db_even.mem_bank[3770],db_odd.mem_bank[3771],db_even.mem_bank[3771],db_odd.mem_bank[3772],db_even.mem_bank[3772],db_odd.mem_bank[3773],db_even.mem_bank[3773],db_odd.mem_bank[3774],db_even.mem_bank[3774],db_odd.mem_bank[3775],db_even.mem_bank[3775],db_odd.mem_bank[3776],db_even.mem_bank[3776],db_odd.mem_bank[3777],db_even.mem_bank[3777],db_odd.mem_bank[3778],db_even.mem_bank[3778],db_odd.mem_bank[3779],db_even.mem_bank[3779],db_odd.mem_bank[3780],db_even.mem_bank[3780],db_odd.mem_bank[3781],db_even.mem_bank[3781],db_odd.mem_bank[3782],db_even.mem_bank[3782],db_odd.mem_bank[3783],db_even.mem_bank[3783],db_odd.mem_bank[3784],db_even.mem_bank[3784],db_odd.mem_bank[3785],db_even.mem_bank[3785],db_odd.mem_bank[3786],db_even.mem_bank[3786],db_odd.mem_bank[3787],db_even.mem_bank[3787],db_odd.mem_bank[3788],db_even.mem_bank[3788],db_odd.mem_bank[3789],db_even.mem_bank[3789],db_odd.mem_bank[3790],db_even.mem_bank[3790],db_odd.mem_bank[3791],db_even.mem_bank[3791],db_odd.mem_bank[3792],db_even.mem_bank[3792],db_odd.mem_bank[3793],db_even.mem_bank[3793],db_odd.mem_bank[3794],db_even.mem_bank[3794],db_odd.mem_bank[3795],db_even.mem_bank[3795],db_odd.mem_bank[3796],db_even.mem_bank[3796],db_odd.mem_bank[3797],db_even.mem_bank[3797],db_odd.mem_bank[3798],db_even.mem_bank[3798],db_odd.mem_bank[3799],db_even.mem_bank[3799],db_odd.mem_bank[3800],db_even.mem_bank[3800],db_odd.mem_bank[3801],db_even.mem_bank[3801],db_odd.mem_bank[3802],db_even.mem_bank[3802],db_odd.mem_bank[3803],db_even.mem_bank[3803],db_odd.mem_bank[3804],db_even.mem_bank[3804],db_odd.mem_bank[3805],db_even.mem_bank[3805],db_odd.mem_bank[3806],db_even.mem_bank[3806],db_odd.mem_bank[3807],db_even.mem_bank[3807],db_odd.mem_bank[3808],db_even.mem_bank[3808],db_odd.mem_bank[3809],db_even.mem_bank[3809],db_odd.mem_bank[3810],db_even.mem_bank[3810],db_odd.mem_bank[3811],db_even.mem_bank[3811],db_odd.mem_bank[3812],db_even.mem_bank[3812],db_odd.mem_bank[3813],db_even.mem_bank[3813],db_odd.mem_bank[3814],db_even.mem_bank[3814],db_odd.mem_bank[3815],db_even.mem_bank[3815],db_odd.mem_bank[3816],db_even.mem_bank[3816],db_odd.mem_bank[3817],db_even.mem_bank[3817],db_odd.mem_bank[3818],db_even.mem_bank[3818],db_odd.mem_bank[3819],db_even.mem_bank[3819],db_odd.mem_bank[3820],db_even.mem_bank[3820],db_odd.mem_bank[3821],db_even.mem_bank[3821],db_odd.mem_bank[3822],db_even.mem_bank[3822],db_odd.mem_bank[3823],db_even.mem_bank[3823],db_odd.mem_bank[3824],db_even.mem_bank[3824],db_odd.mem_bank[3825],db_even.mem_bank[3825],db_odd.mem_bank[3826],db_even.mem_bank[3826],db_odd.mem_bank[3827],db_even.mem_bank[3827],db_odd.mem_bank[3828],db_even.mem_bank[3828],db_odd.mem_bank[3829],db_even.mem_bank[3829],db_odd.mem_bank[3830],db_even.mem_bank[3830],db_odd.mem_bank[3831],db_even.mem_bank[3831],db_odd.mem_bank[3832],db_even.mem_bank[3832],db_odd.mem_bank[3833],db_even.mem_bank[3833],db_odd.mem_bank[3834],db_even.mem_bank[3834],db_odd.mem_bank[3835],db_even.mem_bank[3835],db_odd.mem_bank[3836],db_even.mem_bank[3836],db_odd.mem_bank[3837],db_even.mem_bank[3837],db_odd.mem_bank[3838],db_even.mem_bank[3838],db_odd.mem_bank[3839],db_even.mem_bank[3839],db_odd.mem_bank[3840],db_even.mem_bank[3840],db_odd.mem_bank[3841],db_even.mem_bank[3841],db_odd.mem_bank[3842],db_even.mem_bank[3842],db_odd.mem_bank[3843],db_even.mem_bank[3843],db_odd.mem_bank[3844],db_even.mem_bank[3844],db_odd.mem_bank[3845],db_even.mem_bank[3845],db_odd.mem_bank[3846],db_even.mem_bank[3846],db_odd.mem_bank[3847],db_even.mem_bank[3847],db_odd.mem_bank[3848],db_even.mem_bank[3848],db_odd.mem_bank[3849],db_even.mem_bank[3849],db_odd.mem_bank[3850],db_even.mem_bank[3850],db_odd.mem_bank[3851],db_even.mem_bank[3851],db_odd.mem_bank[3852],db_even.mem_bank[3852],db_odd.mem_bank[3853],db_even.mem_bank[3853],db_odd.mem_bank[3854],db_even.mem_bank[3854],db_odd.mem_bank[3855],db_even.mem_bank[3855],db_odd.mem_bank[3856],db_even.mem_bank[3856],db_odd.mem_bank[3857],db_even.mem_bank[3857],db_odd.mem_bank[3858],db_even.mem_bank[3858],db_odd.mem_bank[3859],db_even.mem_bank[3859],db_odd.mem_bank[3860],db_even.mem_bank[3860],db_odd.mem_bank[3861],db_even.mem_bank[3861],db_odd.mem_bank[3862],db_even.mem_bank[3862],db_odd.mem_bank[3863],db_even.mem_bank[3863],db_odd.mem_bank[3864],db_even.mem_bank[3864],db_odd.mem_bank[3865],db_even.mem_bank[3865],db_odd.mem_bank[3866],db_even.mem_bank[3866],db_odd.mem_bank[3867],db_even.mem_bank[3867],db_odd.mem_bank[3868],db_even.mem_bank[3868],db_odd.mem_bank[3869],db_even.mem_bank[3869],db_odd.mem_bank[3870],db_even.mem_bank[3870],db_odd.mem_bank[3871],db_even.mem_bank[3871],db_odd.mem_bank[3872],db_even.mem_bank[3872],db_odd.mem_bank[3873],db_even.mem_bank[3873],db_odd.mem_bank[3874],db_even.mem_bank[3874],db_odd.mem_bank[3875],db_even.mem_bank[3875],db_odd.mem_bank[3876],db_even.mem_bank[3876],db_odd.mem_bank[3877],db_even.mem_bank[3877],db_odd.mem_bank[3878],db_even.mem_bank[3878],db_odd.mem_bank[3879],db_even.mem_bank[3879],db_odd.mem_bank[3880],db_even.mem_bank[3880],db_odd.mem_bank[3881],db_even.mem_bank[3881],db_odd.mem_bank[3882],db_even.mem_bank[3882],db_odd.mem_bank[3883],db_even.mem_bank[3883],db_odd.mem_bank[3884],db_even.mem_bank[3884],db_odd.mem_bank[3885],db_even.mem_bank[3885],db_odd.mem_bank[3886],db_even.mem_bank[3886],db_odd.mem_bank[3887],db_even.mem_bank[3887],db_odd.mem_bank[3888],db_even.mem_bank[3888],db_odd.mem_bank[3889],db_even.mem_bank[3889],db_odd.mem_bank[3890],db_even.mem_bank[3890],db_odd.mem_bank[3891],db_even.mem_bank[3891],db_odd.mem_bank[3892],db_even.mem_bank[3892],db_odd.mem_bank[3893],db_even.mem_bank[3893],db_odd.mem_bank[3894],db_even.mem_bank[3894],db_odd.mem_bank[3895],db_even.mem_bank[3895],db_odd.mem_bank[3896],db_even.mem_bank[3896],db_odd.mem_bank[3897],db_even.mem_bank[3897],db_odd.mem_bank[3898],db_even.mem_bank[3898],db_odd.mem_bank[3899],db_even.mem_bank[3899],db_odd.mem_bank[3900],db_even.mem_bank[3900],db_odd.mem_bank[3901],db_even.mem_bank[3901],db_odd.mem_bank[3902],db_even.mem_bank[3902],db_odd.mem_bank[3903],db_even.mem_bank[3903],db_odd.mem_bank[3904],db_even.mem_bank[3904],db_odd.mem_bank[3905],db_even.mem_bank[3905],db_odd.mem_bank[3906],db_even.mem_bank[3906],db_odd.mem_bank[3907],db_even.mem_bank[3907],db_odd.mem_bank[3908],db_even.mem_bank[3908],db_odd.mem_bank[3909],db_even.mem_bank[3909],db_odd.mem_bank[3910],db_even.mem_bank[3910],db_odd.mem_bank[3911],db_even.mem_bank[3911],db_odd.mem_bank[3912],db_even.mem_bank[3912],db_odd.mem_bank[3913],db_even.mem_bank[3913],db_odd.mem_bank[3914],db_even.mem_bank[3914],db_odd.mem_bank[3915],db_even.mem_bank[3915],db_odd.mem_bank[3916],db_even.mem_bank[3916],db_odd.mem_bank[3917],db_even.mem_bank[3917],db_odd.mem_bank[3918],db_even.mem_bank[3918],db_odd.mem_bank[3919],db_even.mem_bank[3919],db_odd.mem_bank[3920],db_even.mem_bank[3920],db_odd.mem_bank[3921],db_even.mem_bank[3921],db_odd.mem_bank[3922],db_even.mem_bank[3922],db_odd.mem_bank[3923],db_even.mem_bank[3923],db_odd.mem_bank[3924],db_even.mem_bank[3924],db_odd.mem_bank[3925],db_even.mem_bank[3925],db_odd.mem_bank[3926],db_even.mem_bank[3926],db_odd.mem_bank[3927],db_even.mem_bank[3927],db_odd.mem_bank[3928],db_even.mem_bank[3928],db_odd.mem_bank[3929],db_even.mem_bank[3929],db_odd.mem_bank[3930],db_even.mem_bank[3930],db_odd.mem_bank[3931],db_even.mem_bank[3931],db_odd.mem_bank[3932],db_even.mem_bank[3932],db_odd.mem_bank[3933],db_even.mem_bank[3933],db_odd.mem_bank[3934],db_even.mem_bank[3934],db_odd.mem_bank[3935],db_even.mem_bank[3935],db_odd.mem_bank[3936],db_even.mem_bank[3936],db_odd.mem_bank[3937],db_even.mem_bank[3937],db_odd.mem_bank[3938],db_even.mem_bank[3938],db_odd.mem_bank[3939],db_even.mem_bank[3939],db_odd.mem_bank[3940],db_even.mem_bank[3940],db_odd.mem_bank[3941],db_even.mem_bank[3941],db_odd.mem_bank[3942],db_even.mem_bank[3942],db_odd.mem_bank[3943],db_even.mem_bank[3943],db_odd.mem_bank[3944],db_even.mem_bank[3944],db_odd.mem_bank[3945],db_even.mem_bank[3945],db_odd.mem_bank[3946],db_even.mem_bank[3946],db_odd.mem_bank[3947],db_even.mem_bank[3947],db_odd.mem_bank[3948],db_even.mem_bank[3948],db_odd.mem_bank[3949],db_even.mem_bank[3949],db_odd.mem_bank[3950],db_even.mem_bank[3950],db_odd.mem_bank[3951],db_even.mem_bank[3951],db_odd.mem_bank[3952],db_even.mem_bank[3952],db_odd.mem_bank[3953],db_even.mem_bank[3953],db_odd.mem_bank[3954],db_even.mem_bank[3954],db_odd.mem_bank[3955],db_even.mem_bank[3955],db_odd.mem_bank[3956],db_even.mem_bank[3956],db_odd.mem_bank[3957],db_even.mem_bank[3957],db_odd.mem_bank[3958],db_even.mem_bank[3958],db_odd.mem_bank[3959],db_even.mem_bank[3959],db_odd.mem_bank[3960],db_even.mem_bank[3960],db_odd.mem_bank[3961],db_even.mem_bank[3961],db_odd.mem_bank[3962],db_even.mem_bank[3962],db_odd.mem_bank[3963],db_even.mem_bank[3963],db_odd.mem_bank[3964],db_even.mem_bank[3964],db_odd.mem_bank[3965],db_even.mem_bank[3965],db_odd.mem_bank[3966],db_even.mem_bank[3966],db_odd.mem_bank[3967],db_even.mem_bank[3967],db_odd.mem_bank[3968],db_even.mem_bank[3968],db_odd.mem_bank[3969],db_even.mem_bank[3969],db_odd.mem_bank[3970],db_even.mem_bank[3970],db_odd.mem_bank[3971],db_even.mem_bank[3971],db_odd.mem_bank[3972],db_even.mem_bank[3972],db_odd.mem_bank[3973],db_even.mem_bank[3973],db_odd.mem_bank[3974],db_even.mem_bank[3974],db_odd.mem_bank[3975],db_even.mem_bank[3975],db_odd.mem_bank[3976],db_even.mem_bank[3976],db_odd.mem_bank[3977],db_even.mem_bank[3977],db_odd.mem_bank[3978],db_even.mem_bank[3978],db_odd.mem_bank[3979],db_even.mem_bank[3979],db_odd.mem_bank[3980],db_even.mem_bank[3980],db_odd.mem_bank[3981],db_even.mem_bank[3981],db_odd.mem_bank[3982],db_even.mem_bank[3982],db_odd.mem_bank[3983],db_even.mem_bank[3983],db_odd.mem_bank[3984],db_even.mem_bank[3984],db_odd.mem_bank[3985],db_even.mem_bank[3985],db_odd.mem_bank[3986],db_even.mem_bank[3986],db_odd.mem_bank[3987],db_even.mem_bank[3987],db_odd.mem_bank[3988],db_even.mem_bank[3988],db_odd.mem_bank[3989],db_even.mem_bank[3989],db_odd.mem_bank[3990],db_even.mem_bank[3990],db_odd.mem_bank[3991],db_even.mem_bank[3991],db_odd.mem_bank[3992],db_even.mem_bank[3992],db_odd.mem_bank[3993],db_even.mem_bank[3993],db_odd.mem_bank[3994],db_even.mem_bank[3994],db_odd.mem_bank[3995],db_even.mem_bank[3995],db_odd.mem_bank[3996],db_even.mem_bank[3996],db_odd.mem_bank[3997],db_even.mem_bank[3997],db_odd.mem_bank[3998],db_even.mem_bank[3998],db_odd.mem_bank[3999],db_even.mem_bank[3999],db_odd.mem_bank[4000],db_even.mem_bank[4000],db_odd.mem_bank[4001],db_even.mem_bank[4001],db_odd.mem_bank[4002],db_even.mem_bank[4002],db_odd.mem_bank[4003],db_even.mem_bank[4003],db_odd.mem_bank[4004],db_even.mem_bank[4004],db_odd.mem_bank[4005],db_even.mem_bank[4005],db_odd.mem_bank[4006],db_even.mem_bank[4006],db_odd.mem_bank[4007],db_even.mem_bank[4007],db_odd.mem_bank[4008],db_even.mem_bank[4008],db_odd.mem_bank[4009],db_even.mem_bank[4009],db_odd.mem_bank[4010],db_even.mem_bank[4010],db_odd.mem_bank[4011],db_even.mem_bank[4011],db_odd.mem_bank[4012],db_even.mem_bank[4012],db_odd.mem_bank[4013],db_even.mem_bank[4013],db_odd.mem_bank[4014],db_even.mem_bank[4014],db_odd.mem_bank[4015],db_even.mem_bank[4015],db_odd.mem_bank[4016],db_even.mem_bank[4016],db_odd.mem_bank[4017],db_even.mem_bank[4017],db_odd.mem_bank[4018],db_even.mem_bank[4018],db_odd.mem_bank[4019],db_even.mem_bank[4019],db_odd.mem_bank[4020],db_even.mem_bank[4020],db_odd.mem_bank[4021],db_even.mem_bank[4021],db_odd.mem_bank[4022],db_even.mem_bank[4022],db_odd.mem_bank[4023],db_even.mem_bank[4023],db_odd.mem_bank[4024],db_even.mem_bank[4024],db_odd.mem_bank[4025],db_even.mem_bank[4025],db_odd.mem_bank[4026],db_even.mem_bank[4026],db_odd.mem_bank[4027],db_even.mem_bank[4027],db_odd.mem_bank[4028],db_even.mem_bank[4028],db_odd.mem_bank[4029],db_even.mem_bank[4029],db_odd.mem_bank[4030],db_even.mem_bank[4030],db_odd.mem_bank[4031],db_even.mem_bank[4031],db_odd.mem_bank[4032],db_even.mem_bank[4032],db_odd.mem_bank[4033],db_even.mem_bank[4033],db_odd.mem_bank[4034],db_even.mem_bank[4034],db_odd.mem_bank[4035],db_even.mem_bank[4035],db_odd.mem_bank[4036],db_even.mem_bank[4036],db_odd.mem_bank[4037],db_even.mem_bank[4037],db_odd.mem_bank[4038],db_even.mem_bank[4038],db_odd.mem_bank[4039],db_even.mem_bank[4039],db_odd.mem_bank[4040],db_even.mem_bank[4040],db_odd.mem_bank[4041],db_even.mem_bank[4041],db_odd.mem_bank[4042],db_even.mem_bank[4042],db_odd.mem_bank[4043],db_even.mem_bank[4043],db_odd.mem_bank[4044],db_even.mem_bank[4044],db_odd.mem_bank[4045],db_even.mem_bank[4045],db_odd.mem_bank[4046],db_even.mem_bank[4046],db_odd.mem_bank[4047],db_even.mem_bank[4047],db_odd.mem_bank[4048],db_even.mem_bank[4048],db_odd.mem_bank[4049],db_even.mem_bank[4049],db_odd.mem_bank[4050],db_even.mem_bank[4050],db_odd.mem_bank[4051],db_even.mem_bank[4051],db_odd.mem_bank[4052],db_even.mem_bank[4052],db_odd.mem_bank[4053],db_even.mem_bank[4053],db_odd.mem_bank[4054],db_even.mem_bank[4054],db_odd.mem_bank[4055],db_even.mem_bank[4055],db_odd.mem_bank[4056],db_even.mem_bank[4056],db_odd.mem_bank[4057],db_even.mem_bank[4057],db_odd.mem_bank[4058],db_even.mem_bank[4058],db_odd.mem_bank[4059],db_even.mem_bank[4059],db_odd.mem_bank[4060],db_even.mem_bank[4060],db_odd.mem_bank[4061],db_even.mem_bank[4061],db_odd.mem_bank[4062],db_even.mem_bank[4062],db_odd.mem_bank[4063],db_even.mem_bank[4063],db_odd.mem_bank[4064],db_even.mem_bank[4064],db_odd.mem_bank[4065],db_even.mem_bank[4065],db_odd.mem_bank[4066],db_even.mem_bank[4066],db_odd.mem_bank[4067],db_even.mem_bank[4067],db_odd.mem_bank[4068],db_even.mem_bank[4068],db_odd.mem_bank[4069],db_even.mem_bank[4069],db_odd.mem_bank[4070],db_even.mem_bank[4070],db_odd.mem_bank[4071],db_even.mem_bank[4071],db_odd.mem_bank[4072],db_even.mem_bank[4072],db_odd.mem_bank[4073],db_even.mem_bank[4073],db_odd.mem_bank[4074],db_even.mem_bank[4074],db_odd.mem_bank[4075],db_even.mem_bank[4075],db_odd.mem_bank[4076],db_even.mem_bank[4076],db_odd.mem_bank[4077],db_even.mem_bank[4077],db_odd.mem_bank[4078],db_even.mem_bank[4078],db_odd.mem_bank[4079],db_even.mem_bank[4079],db_odd.mem_bank[4080],db_even.mem_bank[4080],db_odd.mem_bank[4081],db_even.mem_bank[4081],db_odd.mem_bank[4082],db_even.mem_bank[4082],db_odd.mem_bank[4083],db_even.mem_bank[4083],db_odd.mem_bank[4084],db_even.mem_bank[4084],db_odd.mem_bank[4085],db_even.mem_bank[4085],db_odd.mem_bank[4086],db_even.mem_bank[4086],db_odd.mem_bank[4087],db_even.mem_bank[4087],db_odd.mem_bank[4088],db_even.mem_bank[4088],db_odd.mem_bank[4089],db_even.mem_bank[4089],db_odd.mem_bank[4090],db_even.mem_bank[4090],db_odd.mem_bank[4091],db_even.mem_bank[4091],db_odd.mem_bank[4092],db_even.mem_bank[4092],db_odd.mem_bank[4093],db_even.mem_bank[4093],db_odd.mem_bank[4094],db_even.mem_bank[4094],db_odd.mem_bank[4095],db_even.mem_bank[4095]);
  end


endmodule