module d_merge #(
    parameter OOO_TAG_SIZE = 10
    ) (
    
);
    
endmodule