module lsq (

);

endmodule