module ooo_engine_TOP();

endmodule