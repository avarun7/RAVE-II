module regfile_TOP();

endmodule