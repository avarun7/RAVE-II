module dram_top #(parameter CL_SIZE = 128) (
    input clk,
    input rst,

    // I/O FROM INPUT QUEUES
    
    //EVEN SIDE
    //MEM_DATA_Q_in
    input[31:0] addr_in_mem_data_q_even,
    input [CL_SIZE-1:0] data_in_mem_data_q_even,
    input [2:0] operation_in_mem_data_q_even,
    input is_flush_in_mem_data_q_even,
    input alloc_in_mem_data_q_even,
    input [1:0] src_in_mem_data_q_even,
    input [1:0] dest_in_mem_data_q_even,

    output full_out_mem_data_q_even,
    
    //MEM_INSTR_Q_in
    input[31:0] addr_in_mem_instr_q_even,
    input [2:0] operation_in_mem_instr_q_even,
    input is_flush_in_mem_instr_q_even,
    input alloc_in_mem_instr_q_even,
    input [1:0] src_in_mem_instr_q_even,
    input [1:0] dest_in_mem_instr_q_even,

    output full_out_mem_instr_q_even,
    
    //ODD SIDE
    //MEM_DATA_Q_in
    input[31:0] addr_in_mem_data_q_odd,
    input [CL_SIZE-1:0] data_in_mem_data_q_odd,
    input [2:0] operation_in_mem_data_q_odd,
    input is_flush_in_mem_data_q_odd,
    input alloc_in_mem_data_q_odd,
    input [1:0] src_in_mem_data_q_odd,
    input [1:0] dest_in_mem_data_q_odd,

    output full_out_mem_data_q_odd,
    
    //MEM_INSTR_Q_in
    input[31:0] addr_in_mem_instr_q_odd,
    input [2:0] operation_in_mem_instr_q_odd,
    input is_flush_in_mem_instr_q_odd,
    input alloc_in_mem_instr_q_odd,
    input [1:0] src_in_mem_instr_q_odd,
    input [1:0] dest_in_mem_instr_q_odd,

    output full_out_mem_instr_q_odd,

    // I/O to OUTPUT QUEUES

    //EVEN SIDE
    //MEM_DATA_Q_out
    output [31:0] addr_out_mem_data_q_even,
    output [CL_SIZE-1:0] data_out_mem_data_q_even,
    output [2:0] operation_out_mem_data_q_even,
    output is_flush_out_mem_data_q_even,
    output alloc_out_mem_data_q_even,
    output [1:0] src_out_mem_data_q_even,
    output [1:0] dest_out_mem_data_q_even,

    input full_in_mem_data_q_even,

    //ODD SIDE
    //MEM_DATA_Q_out
    output [31:0] addr_out_mem_data_q_odd,
    output  [CL_SIZE-1:0] data_out_mem_data_q_odd,
    output  [2:0] operation_out_mem_data_q_odd,
    output  is_flush_out_mem_data_q_odd,
    output  alloc_out_mem_data_q_odd,
    output  [1:0] src_out_mem_data_q_odd,
    output  [1:0] dest_out_mem_data_q_odd,

    input full_in_mem_data_q_odd
);

       //MEM_DATA_Q_in
wire [31:0] bank_addr_in_mem_data_q_even;
wire  [CL_SIZE-1:0] bank_data_in_mem_data_q_even;
wire  [2:0] bank_operation_in_mem_data_q_even;
wire  bank_is_flush_in_mem_data_q_even;
wire  bank_valid_in_mem_data_q_even;
wire  [1:0] bank_src_in_mem_data_q_even;
wire  [1:0] bank_dest_in_mem_data_q_even;

wire [1:0] dealloc_even, dealloc_odd;
    //MEM_INSTR_Q_in
wire [31:0] bank_addr_in_mem_instr_q_even;
wire  [2:0] bank_operation_in_mem_instr_q_even;
wire  bank_is_flush_in_mem_instr_q_even;
wire  bank_valid_in_mem_instr_q_even;
wire  [1:0] bank_src_in_mem_instr_q_even;
wire  [1:0] bank_dest_in_mem_instr_q_even;
wire [CL_SIZE -1 : 0] bank_data_in_even, bank_data_in_odd;

data_q #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_data_q_even(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_data_q_even),
    .data_in(data_in_mem_data_q_even),
    .operation_in(operation_in_mem_data_q_even),
    .is_flush(is_flush_in_mem_data_q_even),
    .alloc(alloc_in_mem_data_q_even),
    .src(src_in_mem_data_q_even),
    .dest(dest_in_mem_data_q_even),
    //From reciever
    .dealloc(dealloc_even[1]),

    //output sender
    .full(full_out_mem_data_q_even),

    //output reciever
    .addr_out(bank_addr_in_mem_data_q_even),
    .data_out(bank_data_in_mem_data_q_even),
    .operation_out(bank_operation_in_mem_data_q_even),
    .valid(bank_valid_in_mem_data_q_even),
    .src_out(bank_src_in_mem_data_q_even),
    .dest_out(bank_dest_in_mem_data_q_even),
    .is_flush_out(bank_is_flush_in_mem_data_q_even)
);

instr_q  #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_instr_q_even(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_instr_q_even),
    .operation_in(operation_in_mem_instr_q_even),
    .is_flush(is_flush_in_mem_instr_q_even),
    .alloc(alloc_in_mem_instr_q_even),
    .src(src_in_mem_instr_q_even),
    .dest(dest_in_mem_instr_q_even),

    //From reciever
    .dealloc(dealloc_even[0]),

    //output sender
    .full(full_out_mem_instr_q_even),

    //output reciever
    .addr_out(bank_addr_in_mem_instr_q_even),
    .operation_out(bank_operation_in_mem_instr_q_even),
    .valid(bank_valid_in_mem_instr_q_even),
    .src_out(bank_src_in_mem_instr_q_even),
    .dest_out(bank_dest_in_mem_instr_q_even),
    .is_flush_out(bank_is_flush_in_mem_instr_q_even)
);
wire [31:0] bank_addr_in_even;
wire [2:0] bank_operation_in_even;
wire bank_valid_in_even;
// wire [CL_SIZE - 1:0] bank_data_in_even;
wire [1:0] bank_src_in_even;
wire [1:0] bank_dest_in_even;
wire bank_is_flush_in_even;

wire [31:0] bank_addr_in_odd;
wire [2:0] bank_operation_in_odd;
wire bank_valid_in_odd;
// wire [CL_SIZE - 1:0] bank_data_in_odd;
wire [1:0] bank_src_in_odd;
wire [1:0] bank_dest_in_odd;
wire bank_is_flush_in_odd;
queue_arbitrator #(.CL_SIZE(CL_SIZE), .Q_WIDTH(2)) queue_arb_even(
    .addr_in({
        bank_addr_in_mem_data_q_even,
        bank_addr_in_mem_instr_q_even
    }),
    .data_in({
        bank_data_in_mem_data_q_even,
        128'd0
    }),
    .operation_in({
        bank_operation_in_mem_data_q_even,
        bank_operation_in_mem_instr_q_even
    }), 
    .valid_in({
        bank_valid_in_mem_data_q_even,
        bank_valid_in_mem_instr_q_even
    }),
    .src_in({
        bank_src_in_mem_data_q_even,
        bank_src_in_mem_instr_q_even
    }),
    .dest_in({
        bank_dest_in_mem_data_q_even,
        bank_dest_in_mem_instr_q_even
    }),
    .is_flush_in({
        bank_is_flush_in_mem_data_q_even,
        bank_is_flush_in_mem_instr_q_even
    }),
    .stall_in(bank_stall_even),


    .addr_out(      bank_addr_in_even),
    .operation_out( bank_operation_in_even), 
    .valid_out(     bank_valid_in_even),
    .data_out(      bank_data_in_even),
    .src_out(       bank_src_in_even),
    .dest_out(      bank_dest_in_even),
    .is_flush_out(  bank_is_flush_in_even),

    .dealloc(dealloc_even)
);

dram_bank #(.CL_SIZE(CL_SIZE), .file_name(1)) db_even(
.rst(rst),
.clk(clk),

.addr_in(bank_addr_in_even),
.operation_in(bank_operation_in_even),
.valid_in(bank_valid_in_even),
.src_in(bank_src_in_even),
.dest_in(bank_dest_in_even),
.is_flush_in(bank_is_flush_in_even),
.data_in(bank_data_in_even),

.addr_out(addr_out_mem_data_q_even),
.operation_out(operation_out_mem_data_q_even),
.valid_out(alloc_out_mem_data_q_even),
.src_out(src_out_mem_data_q_even),
.dest_out(dest_out_mem_data_q_even),
.is_flush_out(is_flush_out_mem_data_q_even),
.data_out(data_out_mem_data_q_even),

.stall_out(bank_stall_even)
);
      //MEM_DATA_Q_in
wire [31:0] bank_addr_in_mem_data_q_odd;
wire  [CL_SIZE-1:0] bank_data_in_mem_data_q_odd;
wire  [2:0] bank_operation_in_mem_data_q_odd;
wire  bank_is_flush_in_mem_data_q_odd;
wire  bank_valid_in_mem_data_q_odd;
wire  [1:0] bank_src_in_mem_data_q_odd;
wire  [1:0] bank_dest_in_mem_data_q_odd;

    //MEM_INSTR_Q_in
wire [31:0] bank_addr_in_mem_instr_q_odd;
wire  [2:0] bank_operation_in_mem_instr_q_odd;
wire  bank_is_flush_in_mem_instr_q_odd;
wire  bank_valid_in_mem_instr_q_odd;
wire  [1:0] bank_src_in_mem_instr_q_odd;
wire  [1:0] bank_dest_in_mem_instr_q_odd;

data_q #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_data_q_odd(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_data_q_odd),
    .data_in(data_in_mem_data_q_odd),
    .operation_in(operation_in_mem_data_q_odd),
    .is_flush(is_flush_in_mem_data_q_odd),
    .alloc(alloc_in_mem_data_q_odd),
    .src(src_in_mem_data_q_odd),
    .dest(dest_in_mem_data_q_odd),
    //From reciever
    .dealloc(dealloc_odd[1]),

    //output sender
    .full(full_out_mem_data_q_odd),

    //output reciever
    .addr_out(bank_addr_in_mem_data_q_odd),
    .data_out(bank_data_in_mem_data_q_odd),
    .operation_out(bank_operation_in_mem_data_q_odd),
    .valid(bank_valid_in_mem_data_q_odd),
    .src_out(bank_src_in_mem_data_q_odd),
    .dest_out(bank_dest_in_mem_data_q_odd),
    .is_flush_out(bank_is_flush_in_mem_data_q_odd)
);

instr_q  #(.Q_LENGTH(8), .CL_SIZE(CL_SIZE)) mem_instr_q_odd(
    //System     
    .clk(clk),
    .rst(rst),

    //From Sender
    .addr_in(addr_in_mem_instr_q_odd),
    .operation_in(operation_in_mem_instr_q_odd),
    .is_flush(is_flush_in_mem_instr_q_odd),
    .alloc(alloc_in_mem_instr_q_odd),
    .src(src_in_mem_instr_q_odd),
    .dest(dest_in_mem_instr_q_odd),

    //From reciever
    .dealloc(dealloc_odd[0]),

    //output sender
    .full(full_out_mem_instr_q_odd),

    //output reciever
    .addr_out(bank_addr_in_mem_instr_q_odd),
    .operation_out(bank_operation_in_mem_instr_q_odd),
    .valid(bank_valid_in_mem_instr_q_odd),
    .src_out(bank_src_in_mem_instr_q_odd),
    .dest_out(bank_dest_in_mem_instr_q_odd),
    .is_flush_out(bank_is_flush_in_mem_instr_q_odd)
);
queue_arbitrator #(.CL_SIZE(CL_SIZE), .Q_WIDTH(2)) queue_arb_odd(
    .addr_in({
        bank_addr_in_mem_data_q_odd,
        bank_addr_in_mem_instr_q_odd
    }),
    .data_in({
        bank_data_in_mem_data_q_odd,
        128'd0
    }),
    .operation_in({
        bank_operation_in_mem_data_q_odd,
        bank_operation_in_mem_instr_q_odd
    }), 
    .valid_in({
        bank_valid_in_mem_data_q_odd,
        bank_valid_in_mem_instr_q_odd
    }),
    .src_in({
        bank_src_in_mem_data_q_odd,
        bank_src_in_mem_instr_q_odd
    }),
    .dest_in({
        bank_dest_in_mem_data_q_odd,
        bank_dest_in_mem_instr_q_odd
    }),
    .is_flush_in({
        bank_is_flush_in_mem_data_q_odd,
        bank_is_flush_in_mem_instr_q_odd
    }),

    .stall_in(bank_stall_odd),

    .addr_out(bank_addr_in_odd),
    .operation_out(bank_operation_in_odd), 
    .valid_out(bank_valid_in_odd),
    .data_out(bank_data_in_odd),
    .src_out(bank_src_in_odd),
    .dest_out(bank_dest_in_odd),
    .is_flush_out(bank_is_flush_in_odd),

    .dealloc(dealloc_odd)
);

dram_bank #(.CL_SIZE(128), .file_name(2)) db_odd(
.rst(rst),
.clk(clk),

.addr_in(bank_addr_in_odd),
.operation_in(bank_operation_in_odd),
.valid_in(bank_valid_in_odd),
.src_in(bank_src_in_odd),
.dest_in(bank_dest_in_odd),
.is_flush_in(bank_is_flush_in_odd),
.data_in(bank_data_in_odd),

.addr_out(addr_out_mem_data_q_odd),
.operation_out(operation_out_mem_data_q_odd),
.valid_out(alloc_out_mem_data_q_odd),
.src_out(src_out_mem_data_q_odd),
.dest_out(dest_out_mem_data_q_odd),
.is_flush_out(is_flush_out_mem_data_q_odd),
.data_out(data_out_mem_data_q_odd),

.stall_out(bank_stall_odd)
);


integer file;
  integer count = 0;
initial begin
    file = $fopen("out/MEM_FINAL.csv", "w");
    if (file == 0) begin
      $display("Error: Unable to open file.");
      $stop;
    end
    $fdisplay(file, "Little Endian - Smallest address on the right, largest address left\n");

    #400
    $fdisplay(file, "0x0,0x%h_0x%h", db_odd.mem_bank[0],db_even.mem_bank[0]);
$fdisplay(file, "0x20,0x%h_0x%h", db_odd.mem_bank[1],db_even.mem_bank[1]);
$fdisplay(file, "0x40,0x%h_0x%h", db_odd.mem_bank[2],db_even.mem_bank[2]);
$fdisplay(file, "0x60,0x%h_0x%h", db_odd.mem_bank[3],db_even.mem_bank[3]);
$fdisplay(file, "0x80,0x%h_0x%h", db_odd.mem_bank[4],db_even.mem_bank[4]);
$fdisplay(file, "0xA0,0x%h_0x%h", db_odd.mem_bank[5],db_even.mem_bank[5]);
$fdisplay(file, "0xC0,0x%h_0x%h", db_odd.mem_bank[6],db_even.mem_bank[6]);
$fdisplay(file, "0xE0,0x%h_0x%h", db_odd.mem_bank[7],db_even.mem_bank[7]);
$fdisplay(file, "0x100,0x%h_0x%h", db_odd.mem_bank[8],db_even.mem_bank[8]);
$fdisplay(file, "0x120,0x%h_0x%h", db_odd.mem_bank[9],db_even.mem_bank[9]);
$fdisplay(file, "0x140,0x%h_0x%h", db_odd.mem_bank[10],db_even.mem_bank[10]);
$fdisplay(file, "0x160,0x%h_0x%h", db_odd.mem_bank[11],db_even.mem_bank[11]);
$fdisplay(file, "0x180,0x%h_0x%h", db_odd.mem_bank[12],db_even.mem_bank[12]);
$fdisplay(file, "0x1A0,0x%h_0x%h", db_odd.mem_bank[13],db_even.mem_bank[13]);
$fdisplay(file, "0x1C0,0x%h_0x%h", db_odd.mem_bank[14],db_even.mem_bank[14]);
$fdisplay(file, "0x1E0,0x%h_0x%h", db_odd.mem_bank[15],db_even.mem_bank[15]);
$fdisplay(file, "0x200,0x%h_0x%h", db_odd.mem_bank[16],db_even.mem_bank[16]);
$fdisplay(file, "0x220,0x%h_0x%h", db_odd.mem_bank[17],db_even.mem_bank[17]);
$fdisplay(file, "0x240,0x%h_0x%h", db_odd.mem_bank[18],db_even.mem_bank[18]);
$fdisplay(file, "0x260,0x%h_0x%h", db_odd.mem_bank[19],db_even.mem_bank[19]);
$fdisplay(file, "0x280,0x%h_0x%h", db_odd.mem_bank[20],db_even.mem_bank[20]);
$fdisplay(file, "0x2A0,0x%h_0x%h", db_odd.mem_bank[21],db_even.mem_bank[21]);
$fdisplay(file, "0x2C0,0x%h_0x%h", db_odd.mem_bank[22],db_even.mem_bank[22]);
$fdisplay(file, "0x2E0,0x%h_0x%h", db_odd.mem_bank[23],db_even.mem_bank[23]);
$fdisplay(file, "0x300,0x%h_0x%h", db_odd.mem_bank[24],db_even.mem_bank[24]);
$fdisplay(file, "0x320,0x%h_0x%h", db_odd.mem_bank[25],db_even.mem_bank[25]);
$fdisplay(file, "0x340,0x%h_0x%h", db_odd.mem_bank[26],db_even.mem_bank[26]);
$fdisplay(file, "0x360,0x%h_0x%h", db_odd.mem_bank[27],db_even.mem_bank[27]);
$fdisplay(file, "0x380,0x%h_0x%h", db_odd.mem_bank[28],db_even.mem_bank[28]);
$fdisplay(file, "0x3A0,0x%h_0x%h", db_odd.mem_bank[29],db_even.mem_bank[29]);
$fdisplay(file, "0x3C0,0x%h_0x%h", db_odd.mem_bank[30],db_even.mem_bank[30]);
$fdisplay(file, "0x3E0,0x%h_0x%h", db_odd.mem_bank[31],db_even.mem_bank[31]);
$fdisplay(file, "0x400,0x%h_0x%h", db_odd.mem_bank[32],db_even.mem_bank[32]);
$fdisplay(file, "0x420,0x%h_0x%h", db_odd.mem_bank[33],db_even.mem_bank[33]);
$fdisplay(file, "0x440,0x%h_0x%h", db_odd.mem_bank[34],db_even.mem_bank[34]);
$fdisplay(file, "0x460,0x%h_0x%h", db_odd.mem_bank[35],db_even.mem_bank[35]);
$fdisplay(file, "0x480,0x%h_0x%h", db_odd.mem_bank[36],db_even.mem_bank[36]);
$fdisplay(file, "0x4A0,0x%h_0x%h", db_odd.mem_bank[37],db_even.mem_bank[37]);
$fdisplay(file, "0x4C0,0x%h_0x%h", db_odd.mem_bank[38],db_even.mem_bank[38]);
$fdisplay(file, "0x4E0,0x%h_0x%h", db_odd.mem_bank[39],db_even.mem_bank[39]);
$fdisplay(file, "0x500,0x%h_0x%h", db_odd.mem_bank[40],db_even.mem_bank[40]);
$fdisplay(file, "0x520,0x%h_0x%h", db_odd.mem_bank[41],db_even.mem_bank[41]);
$fdisplay(file, "0x540,0x%h_0x%h", db_odd.mem_bank[42],db_even.mem_bank[42]);
$fdisplay(file, "0x560,0x%h_0x%h", db_odd.mem_bank[43],db_even.mem_bank[43]);
$fdisplay(file, "0x580,0x%h_0x%h", db_odd.mem_bank[44],db_even.mem_bank[44]);
$fdisplay(file, "0x5A0,0x%h_0x%h", db_odd.mem_bank[45],db_even.mem_bank[45]);
$fdisplay(file, "0x5C0,0x%h_0x%h", db_odd.mem_bank[46],db_even.mem_bank[46]);
$fdisplay(file, "0x5E0,0x%h_0x%h", db_odd.mem_bank[47],db_even.mem_bank[47]);
$fdisplay(file, "0x600,0x%h_0x%h", db_odd.mem_bank[48],db_even.mem_bank[48]);
$fdisplay(file, "0x620,0x%h_0x%h", db_odd.mem_bank[49],db_even.mem_bank[49]);
$fdisplay(file, "0x640,0x%h_0x%h", db_odd.mem_bank[50],db_even.mem_bank[50]);
$fdisplay(file, "0x660,0x%h_0x%h", db_odd.mem_bank[51],db_even.mem_bank[51]);
$fdisplay(file, "0x680,0x%h_0x%h", db_odd.mem_bank[52],db_even.mem_bank[52]);
$fdisplay(file, "0x6A0,0x%h_0x%h", db_odd.mem_bank[53],db_even.mem_bank[53]);
$fdisplay(file, "0x6C0,0x%h_0x%h", db_odd.mem_bank[54],db_even.mem_bank[54]);
$fdisplay(file, "0x6E0,0x%h_0x%h", db_odd.mem_bank[55],db_even.mem_bank[55]);
$fdisplay(file, "0x700,0x%h_0x%h", db_odd.mem_bank[56],db_even.mem_bank[56]);
$fdisplay(file, "0x720,0x%h_0x%h", db_odd.mem_bank[57],db_even.mem_bank[57]);
$fdisplay(file, "0x740,0x%h_0x%h", db_odd.mem_bank[58],db_even.mem_bank[58]);
$fdisplay(file, "0x760,0x%h_0x%h", db_odd.mem_bank[59],db_even.mem_bank[59]);
$fdisplay(file, "0x780,0x%h_0x%h", db_odd.mem_bank[60],db_even.mem_bank[60]);
$fdisplay(file, "0x7A0,0x%h_0x%h", db_odd.mem_bank[61],db_even.mem_bank[61]);
$fdisplay(file, "0x7C0,0x%h_0x%h", db_odd.mem_bank[62],db_even.mem_bank[62]);
$fdisplay(file, "0x7E0,0x%h_0x%h", db_odd.mem_bank[63],db_even.mem_bank[63]);
$fdisplay(file, "0x800,0x%h_0x%h", db_odd.mem_bank[64],db_even.mem_bank[64]);
$fdisplay(file, "0x820,0x%h_0x%h", db_odd.mem_bank[65],db_even.mem_bank[65]);
$fdisplay(file, "0x840,0x%h_0x%h", db_odd.mem_bank[66],db_even.mem_bank[66]);
$fdisplay(file, "0x860,0x%h_0x%h", db_odd.mem_bank[67],db_even.mem_bank[67]);
$fdisplay(file, "0x880,0x%h_0x%h", db_odd.mem_bank[68],db_even.mem_bank[68]);
$fdisplay(file, "0x8A0,0x%h_0x%h", db_odd.mem_bank[69],db_even.mem_bank[69]);
$fdisplay(file, "0x8C0,0x%h_0x%h", db_odd.mem_bank[70],db_even.mem_bank[70]);
$fdisplay(file, "0x8E0,0x%h_0x%h", db_odd.mem_bank[71],db_even.mem_bank[71]);
$fdisplay(file, "0x900,0x%h_0x%h", db_odd.mem_bank[72],db_even.mem_bank[72]);
$fdisplay(file, "0x920,0x%h_0x%h", db_odd.mem_bank[73],db_even.mem_bank[73]);
$fdisplay(file, "0x940,0x%h_0x%h", db_odd.mem_bank[74],db_even.mem_bank[74]);
$fdisplay(file, "0x960,0x%h_0x%h", db_odd.mem_bank[75],db_even.mem_bank[75]);
$fdisplay(file, "0x980,0x%h_0x%h", db_odd.mem_bank[76],db_even.mem_bank[76]);
$fdisplay(file, "0x9A0,0x%h_0x%h", db_odd.mem_bank[77],db_even.mem_bank[77]);
$fdisplay(file, "0x9C0,0x%h_0x%h", db_odd.mem_bank[78],db_even.mem_bank[78]);
$fdisplay(file, "0x9E0,0x%h_0x%h", db_odd.mem_bank[79],db_even.mem_bank[79]);
$fdisplay(file, "0xA00,0x%h_0x%h", db_odd.mem_bank[80],db_even.mem_bank[80]);
$fdisplay(file, "0xA20,0x%h_0x%h", db_odd.mem_bank[81],db_even.mem_bank[81]);
$fdisplay(file, "0xA40,0x%h_0x%h", db_odd.mem_bank[82],db_even.mem_bank[82]);
$fdisplay(file, "0xA60,0x%h_0x%h", db_odd.mem_bank[83],db_even.mem_bank[83]);
$fdisplay(file, "0xA80,0x%h_0x%h", db_odd.mem_bank[84],db_even.mem_bank[84]);
$fdisplay(file, "0xAA0,0x%h_0x%h", db_odd.mem_bank[85],db_even.mem_bank[85]);
$fdisplay(file, "0xAC0,0x%h_0x%h", db_odd.mem_bank[86],db_even.mem_bank[86]);
$fdisplay(file, "0xAE0,0x%h_0x%h", db_odd.mem_bank[87],db_even.mem_bank[87]);
$fdisplay(file, "0xB00,0x%h_0x%h", db_odd.mem_bank[88],db_even.mem_bank[88]);
$fdisplay(file, "0xB20,0x%h_0x%h", db_odd.mem_bank[89],db_even.mem_bank[89]);
$fdisplay(file, "0xB40,0x%h_0x%h", db_odd.mem_bank[90],db_even.mem_bank[90]);
$fdisplay(file, "0xB60,0x%h_0x%h", db_odd.mem_bank[91],db_even.mem_bank[91]);
$fdisplay(file, "0xB80,0x%h_0x%h", db_odd.mem_bank[92],db_even.mem_bank[92]);
$fdisplay(file, "0xBA0,0x%h_0x%h", db_odd.mem_bank[93],db_even.mem_bank[93]);
$fdisplay(file, "0xBC0,0x%h_0x%h", db_odd.mem_bank[94],db_even.mem_bank[94]);
$fdisplay(file, "0xBE0,0x%h_0x%h", db_odd.mem_bank[95],db_even.mem_bank[95]);
$fdisplay(file, "0xC00,0x%h_0x%h", db_odd.mem_bank[96],db_even.mem_bank[96]);
$fdisplay(file, "0xC20,0x%h_0x%h", db_odd.mem_bank[97],db_even.mem_bank[97]);
$fdisplay(file, "0xC40,0x%h_0x%h", db_odd.mem_bank[98],db_even.mem_bank[98]);
$fdisplay(file, "0xC60,0x%h_0x%h", db_odd.mem_bank[99],db_even.mem_bank[99]);
$fdisplay(file, "0xC80,0x%h_0x%h", db_odd.mem_bank[100],db_even.mem_bank[100]);
$fdisplay(file, "0xCA0,0x%h_0x%h", db_odd.mem_bank[101],db_even.mem_bank[101]);
$fdisplay(file, "0xCC0,0x%h_0x%h", db_odd.mem_bank[102],db_even.mem_bank[102]);
$fdisplay(file, "0xCE0,0x%h_0x%h", db_odd.mem_bank[103],db_even.mem_bank[103]);
$fdisplay(file, "0xD00,0x%h_0x%h", db_odd.mem_bank[104],db_even.mem_bank[104]);
$fdisplay(file, "0xD20,0x%h_0x%h", db_odd.mem_bank[105],db_even.mem_bank[105]);
$fdisplay(file, "0xD40,0x%h_0x%h", db_odd.mem_bank[106],db_even.mem_bank[106]);
$fdisplay(file, "0xD60,0x%h_0x%h", db_odd.mem_bank[107],db_even.mem_bank[107]);
$fdisplay(file, "0xD80,0x%h_0x%h", db_odd.mem_bank[108],db_even.mem_bank[108]);
$fdisplay(file, "0xDA0,0x%h_0x%h", db_odd.mem_bank[109],db_even.mem_bank[109]);
$fdisplay(file, "0xDC0,0x%h_0x%h", db_odd.mem_bank[110],db_even.mem_bank[110]);
$fdisplay(file, "0xDE0,0x%h_0x%h", db_odd.mem_bank[111],db_even.mem_bank[111]);
$fdisplay(file, "0xE00,0x%h_0x%h", db_odd.mem_bank[112],db_even.mem_bank[112]);
$fdisplay(file, "0xE20,0x%h_0x%h", db_odd.mem_bank[113],db_even.mem_bank[113]);
$fdisplay(file, "0xE40,0x%h_0x%h", db_odd.mem_bank[114],db_even.mem_bank[114]);
$fdisplay(file, "0xE60,0x%h_0x%h", db_odd.mem_bank[115],db_even.mem_bank[115]);
$fdisplay(file, "0xE80,0x%h_0x%h", db_odd.mem_bank[116],db_even.mem_bank[116]);
$fdisplay(file, "0xEA0,0x%h_0x%h", db_odd.mem_bank[117],db_even.mem_bank[117]);
$fdisplay(file, "0xEC0,0x%h_0x%h", db_odd.mem_bank[118],db_even.mem_bank[118]);
$fdisplay(file, "0xEE0,0x%h_0x%h", db_odd.mem_bank[119],db_even.mem_bank[119]);
$fdisplay(file, "0xF00,0x%h_0x%h", db_odd.mem_bank[120],db_even.mem_bank[120]);
$fdisplay(file, "0xF20,0x%h_0x%h", db_odd.mem_bank[121],db_even.mem_bank[121]);
$fdisplay(file, "0xF40,0x%h_0x%h", db_odd.mem_bank[122],db_even.mem_bank[122]);
$fdisplay(file, "0xF60,0x%h_0x%h", db_odd.mem_bank[123],db_even.mem_bank[123]);
$fdisplay(file, "0xF80,0x%h_0x%h", db_odd.mem_bank[124],db_even.mem_bank[124]);
$fdisplay(file, "0xFA0,0x%h_0x%h", db_odd.mem_bank[125],db_even.mem_bank[125]);
$fdisplay(file, "0xFC0,0x%h_0x%h", db_odd.mem_bank[126],db_even.mem_bank[126]);
$fdisplay(file, "0xFE0,0x%h_0x%h", db_odd.mem_bank[127],db_even.mem_bank[127]);
$fdisplay(file, "0x1000,0x%h_0x%h", db_odd.mem_bank[128],db_even.mem_bank[128]);
$fdisplay(file, "0x1020,0x%h_0x%h", db_odd.mem_bank[129],db_even.mem_bank[129]);
$fdisplay(file, "0x1040,0x%h_0x%h", db_odd.mem_bank[130],db_even.mem_bank[130]);
$fdisplay(file, "0x1060,0x%h_0x%h", db_odd.mem_bank[131],db_even.mem_bank[131]);
$fdisplay(file, "0x1080,0x%h_0x%h", db_odd.mem_bank[132],db_even.mem_bank[132]);
$fdisplay(file, "0x10A0,0x%h_0x%h", db_odd.mem_bank[133],db_even.mem_bank[133]);
$fdisplay(file, "0x10C0,0x%h_0x%h", db_odd.mem_bank[134],db_even.mem_bank[134]);
$fdisplay(file, "0x10E0,0x%h_0x%h", db_odd.mem_bank[135],db_even.mem_bank[135]);
$fdisplay(file, "0x1100,0x%h_0x%h", db_odd.mem_bank[136],db_even.mem_bank[136]);
$fdisplay(file, "0x1120,0x%h_0x%h", db_odd.mem_bank[137],db_even.mem_bank[137]);
$fdisplay(file, "0x1140,0x%h_0x%h", db_odd.mem_bank[138],db_even.mem_bank[138]);
$fdisplay(file, "0x1160,0x%h_0x%h", db_odd.mem_bank[139],db_even.mem_bank[139]);
$fdisplay(file, "0x1180,0x%h_0x%h", db_odd.mem_bank[140],db_even.mem_bank[140]);
$fdisplay(file, "0x11A0,0x%h_0x%h", db_odd.mem_bank[141],db_even.mem_bank[141]);
$fdisplay(file, "0x11C0,0x%h_0x%h", db_odd.mem_bank[142],db_even.mem_bank[142]);
$fdisplay(file, "0x11E0,0x%h_0x%h", db_odd.mem_bank[143],db_even.mem_bank[143]);
$fdisplay(file, "0x1200,0x%h_0x%h", db_odd.mem_bank[144],db_even.mem_bank[144]);
$fdisplay(file, "0x1220,0x%h_0x%h", db_odd.mem_bank[145],db_even.mem_bank[145]);
$fdisplay(file, "0x1240,0x%h_0x%h", db_odd.mem_bank[146],db_even.mem_bank[146]);
$fdisplay(file, "0x1260,0x%h_0x%h", db_odd.mem_bank[147],db_even.mem_bank[147]);
$fdisplay(file, "0x1280,0x%h_0x%h", db_odd.mem_bank[148],db_even.mem_bank[148]);
$fdisplay(file, "0x12A0,0x%h_0x%h", db_odd.mem_bank[149],db_even.mem_bank[149]);
$fdisplay(file, "0x12C0,0x%h_0x%h", db_odd.mem_bank[150],db_even.mem_bank[150]);
$fdisplay(file, "0x12E0,0x%h_0x%h", db_odd.mem_bank[151],db_even.mem_bank[151]);
$fdisplay(file, "0x1300,0x%h_0x%h", db_odd.mem_bank[152],db_even.mem_bank[152]);
$fdisplay(file, "0x1320,0x%h_0x%h", db_odd.mem_bank[153],db_even.mem_bank[153]);
$fdisplay(file, "0x1340,0x%h_0x%h", db_odd.mem_bank[154],db_even.mem_bank[154]);
$fdisplay(file, "0x1360,0x%h_0x%h", db_odd.mem_bank[155],db_even.mem_bank[155]);
$fdisplay(file, "0x1380,0x%h_0x%h", db_odd.mem_bank[156],db_even.mem_bank[156]);
$fdisplay(file, "0x13A0,0x%h_0x%h", db_odd.mem_bank[157],db_even.mem_bank[157]);
$fdisplay(file, "0x13C0,0x%h_0x%h", db_odd.mem_bank[158],db_even.mem_bank[158]);
$fdisplay(file, "0x13E0,0x%h_0x%h", db_odd.mem_bank[159],db_even.mem_bank[159]);
$fdisplay(file, "0x1400,0x%h_0x%h", db_odd.mem_bank[160],db_even.mem_bank[160]);
$fdisplay(file, "0x1420,0x%h_0x%h", db_odd.mem_bank[161],db_even.mem_bank[161]);
$fdisplay(file, "0x1440,0x%h_0x%h", db_odd.mem_bank[162],db_even.mem_bank[162]);
$fdisplay(file, "0x1460,0x%h_0x%h", db_odd.mem_bank[163],db_even.mem_bank[163]);
$fdisplay(file, "0x1480,0x%h_0x%h", db_odd.mem_bank[164],db_even.mem_bank[164]);
$fdisplay(file, "0x14A0,0x%h_0x%h", db_odd.mem_bank[165],db_even.mem_bank[165]);
$fdisplay(file, "0x14C0,0x%h_0x%h", db_odd.mem_bank[166],db_even.mem_bank[166]);
$fdisplay(file, "0x14E0,0x%h_0x%h", db_odd.mem_bank[167],db_even.mem_bank[167]);
$fdisplay(file, "0x1500,0x%h_0x%h", db_odd.mem_bank[168],db_even.mem_bank[168]);
$fdisplay(file, "0x1520,0x%h_0x%h", db_odd.mem_bank[169],db_even.mem_bank[169]);
$fdisplay(file, "0x1540,0x%h_0x%h", db_odd.mem_bank[170],db_even.mem_bank[170]);
$fdisplay(file, "0x1560,0x%h_0x%h", db_odd.mem_bank[171],db_even.mem_bank[171]);
$fdisplay(file, "0x1580,0x%h_0x%h", db_odd.mem_bank[172],db_even.mem_bank[172]);
$fdisplay(file, "0x15A0,0x%h_0x%h", db_odd.mem_bank[173],db_even.mem_bank[173]);
$fdisplay(file, "0x15C0,0x%h_0x%h", db_odd.mem_bank[174],db_even.mem_bank[174]);
$fdisplay(file, "0x15E0,0x%h_0x%h", db_odd.mem_bank[175],db_even.mem_bank[175]);
$fdisplay(file, "0x1600,0x%h_0x%h", db_odd.mem_bank[176],db_even.mem_bank[176]);
$fdisplay(file, "0x1620,0x%h_0x%h", db_odd.mem_bank[177],db_even.mem_bank[177]);
$fdisplay(file, "0x1640,0x%h_0x%h", db_odd.mem_bank[178],db_even.mem_bank[178]);
$fdisplay(file, "0x1660,0x%h_0x%h", db_odd.mem_bank[179],db_even.mem_bank[179]);
$fdisplay(file, "0x1680,0x%h_0x%h", db_odd.mem_bank[180],db_even.mem_bank[180]);
$fdisplay(file, "0x16A0,0x%h_0x%h", db_odd.mem_bank[181],db_even.mem_bank[181]);
$fdisplay(file, "0x16C0,0x%h_0x%h", db_odd.mem_bank[182],db_even.mem_bank[182]);
$fdisplay(file, "0x16E0,0x%h_0x%h", db_odd.mem_bank[183],db_even.mem_bank[183]);
$fdisplay(file, "0x1700,0x%h_0x%h", db_odd.mem_bank[184],db_even.mem_bank[184]);
$fdisplay(file, "0x1720,0x%h_0x%h", db_odd.mem_bank[185],db_even.mem_bank[185]);
$fdisplay(file, "0x1740,0x%h_0x%h", db_odd.mem_bank[186],db_even.mem_bank[186]);
$fdisplay(file, "0x1760,0x%h_0x%h", db_odd.mem_bank[187],db_even.mem_bank[187]);
$fdisplay(file, "0x1780,0x%h_0x%h", db_odd.mem_bank[188],db_even.mem_bank[188]);
$fdisplay(file, "0x17A0,0x%h_0x%h", db_odd.mem_bank[189],db_even.mem_bank[189]);
$fdisplay(file, "0x17C0,0x%h_0x%h", db_odd.mem_bank[190],db_even.mem_bank[190]);
$fdisplay(file, "0x17E0,0x%h_0x%h", db_odd.mem_bank[191],db_even.mem_bank[191]);
$fdisplay(file, "0x1800,0x%h_0x%h", db_odd.mem_bank[192],db_even.mem_bank[192]);
$fdisplay(file, "0x1820,0x%h_0x%h", db_odd.mem_bank[193],db_even.mem_bank[193]);
$fdisplay(file, "0x1840,0x%h_0x%h", db_odd.mem_bank[194],db_even.mem_bank[194]);
$fdisplay(file, "0x1860,0x%h_0x%h", db_odd.mem_bank[195],db_even.mem_bank[195]);
$fdisplay(file, "0x1880,0x%h_0x%h", db_odd.mem_bank[196],db_even.mem_bank[196]);
$fdisplay(file, "0x18A0,0x%h_0x%h", db_odd.mem_bank[197],db_even.mem_bank[197]);
$fdisplay(file, "0x18C0,0x%h_0x%h", db_odd.mem_bank[198],db_even.mem_bank[198]);
$fdisplay(file, "0x18E0,0x%h_0x%h", db_odd.mem_bank[199],db_even.mem_bank[199]);
$fdisplay(file, "0x1900,0x%h_0x%h", db_odd.mem_bank[200],db_even.mem_bank[200]);
$fdisplay(file, "0x1920,0x%h_0x%h", db_odd.mem_bank[201],db_even.mem_bank[201]);
$fdisplay(file, "0x1940,0x%h_0x%h", db_odd.mem_bank[202],db_even.mem_bank[202]);
$fdisplay(file, "0x1960,0x%h_0x%h", db_odd.mem_bank[203],db_even.mem_bank[203]);
$fdisplay(file, "0x1980,0x%h_0x%h", db_odd.mem_bank[204],db_even.mem_bank[204]);
$fdisplay(file, "0x19A0,0x%h_0x%h", db_odd.mem_bank[205],db_even.mem_bank[205]);
$fdisplay(file, "0x19C0,0x%h_0x%h", db_odd.mem_bank[206],db_even.mem_bank[206]);
$fdisplay(file, "0x19E0,0x%h_0x%h", db_odd.mem_bank[207],db_even.mem_bank[207]);
$fdisplay(file, "0x1A00,0x%h_0x%h", db_odd.mem_bank[208],db_even.mem_bank[208]);
$fdisplay(file, "0x1A20,0x%h_0x%h", db_odd.mem_bank[209],db_even.mem_bank[209]);
$fdisplay(file, "0x1A40,0x%h_0x%h", db_odd.mem_bank[210],db_even.mem_bank[210]);
$fdisplay(file, "0x1A60,0x%h_0x%h", db_odd.mem_bank[211],db_even.mem_bank[211]);
$fdisplay(file, "0x1A80,0x%h_0x%h", db_odd.mem_bank[212],db_even.mem_bank[212]);
$fdisplay(file, "0x1AA0,0x%h_0x%h", db_odd.mem_bank[213],db_even.mem_bank[213]);
$fdisplay(file, "0x1AC0,0x%h_0x%h", db_odd.mem_bank[214],db_even.mem_bank[214]);
$fdisplay(file, "0x1AE0,0x%h_0x%h", db_odd.mem_bank[215],db_even.mem_bank[215]);
$fdisplay(file, "0x1B00,0x%h_0x%h", db_odd.mem_bank[216],db_even.mem_bank[216]);
$fdisplay(file, "0x1B20,0x%h_0x%h", db_odd.mem_bank[217],db_even.mem_bank[217]);
$fdisplay(file, "0x1B40,0x%h_0x%h", db_odd.mem_bank[218],db_even.mem_bank[218]);
$fdisplay(file, "0x1B60,0x%h_0x%h", db_odd.mem_bank[219],db_even.mem_bank[219]);
$fdisplay(file, "0x1B80,0x%h_0x%h", db_odd.mem_bank[220],db_even.mem_bank[220]);
$fdisplay(file, "0x1BA0,0x%h_0x%h", db_odd.mem_bank[221],db_even.mem_bank[221]);
$fdisplay(file, "0x1BC0,0x%h_0x%h", db_odd.mem_bank[222],db_even.mem_bank[222]);
$fdisplay(file, "0x1BE0,0x%h_0x%h", db_odd.mem_bank[223],db_even.mem_bank[223]);
$fdisplay(file, "0x1C00,0x%h_0x%h", db_odd.mem_bank[224],db_even.mem_bank[224]);
$fdisplay(file, "0x1C20,0x%h_0x%h", db_odd.mem_bank[225],db_even.mem_bank[225]);
$fdisplay(file, "0x1C40,0x%h_0x%h", db_odd.mem_bank[226],db_even.mem_bank[226]);
$fdisplay(file, "0x1C60,0x%h_0x%h", db_odd.mem_bank[227],db_even.mem_bank[227]);
$fdisplay(file, "0x1C80,0x%h_0x%h", db_odd.mem_bank[228],db_even.mem_bank[228]);
$fdisplay(file, "0x1CA0,0x%h_0x%h", db_odd.mem_bank[229],db_even.mem_bank[229]);
$fdisplay(file, "0x1CC0,0x%h_0x%h", db_odd.mem_bank[230],db_even.mem_bank[230]);
$fdisplay(file, "0x1CE0,0x%h_0x%h", db_odd.mem_bank[231],db_even.mem_bank[231]);
$fdisplay(file, "0x1D00,0x%h_0x%h", db_odd.mem_bank[232],db_even.mem_bank[232]);
$fdisplay(file, "0x1D20,0x%h_0x%h", db_odd.mem_bank[233],db_even.mem_bank[233]);
$fdisplay(file, "0x1D40,0x%h_0x%h", db_odd.mem_bank[234],db_even.mem_bank[234]);
$fdisplay(file, "0x1D60,0x%h_0x%h", db_odd.mem_bank[235],db_even.mem_bank[235]);
$fdisplay(file, "0x1D80,0x%h_0x%h", db_odd.mem_bank[236],db_even.mem_bank[236]);
$fdisplay(file, "0x1DA0,0x%h_0x%h", db_odd.mem_bank[237],db_even.mem_bank[237]);
$fdisplay(file, "0x1DC0,0x%h_0x%h", db_odd.mem_bank[238],db_even.mem_bank[238]);
$fdisplay(file, "0x1DE0,0x%h_0x%h", db_odd.mem_bank[239],db_even.mem_bank[239]);
$fdisplay(file, "0x1E00,0x%h_0x%h", db_odd.mem_bank[240],db_even.mem_bank[240]);
$fdisplay(file, "0x1E20,0x%h_0x%h", db_odd.mem_bank[241],db_even.mem_bank[241]);
$fdisplay(file, "0x1E40,0x%h_0x%h", db_odd.mem_bank[242],db_even.mem_bank[242]);
$fdisplay(file, "0x1E60,0x%h_0x%h", db_odd.mem_bank[243],db_even.mem_bank[243]);
$fdisplay(file, "0x1E80,0x%h_0x%h", db_odd.mem_bank[244],db_even.mem_bank[244]);
$fdisplay(file, "0x1EA0,0x%h_0x%h", db_odd.mem_bank[245],db_even.mem_bank[245]);
$fdisplay(file, "0x1EC0,0x%h_0x%h", db_odd.mem_bank[246],db_even.mem_bank[246]);
$fdisplay(file, "0x1EE0,0x%h_0x%h", db_odd.mem_bank[247],db_even.mem_bank[247]);
$fdisplay(file, "0x1F00,0x%h_0x%h", db_odd.mem_bank[248],db_even.mem_bank[248]);
$fdisplay(file, "0x1F20,0x%h_0x%h", db_odd.mem_bank[249],db_even.mem_bank[249]);
$fdisplay(file, "0x1F40,0x%h_0x%h", db_odd.mem_bank[250],db_even.mem_bank[250]);
$fdisplay(file, "0x1F60,0x%h_0x%h", db_odd.mem_bank[251],db_even.mem_bank[251]);
$fdisplay(file, "0x1F80,0x%h_0x%h", db_odd.mem_bank[252],db_even.mem_bank[252]);
$fdisplay(file, "0x1FA0,0x%h_0x%h", db_odd.mem_bank[253],db_even.mem_bank[253]);
$fdisplay(file, "0x1FC0,0x%h_0x%h", db_odd.mem_bank[254],db_even.mem_bank[254]);
$fdisplay(file, "0x1FE0,0x%h_0x%h", db_odd.mem_bank[255],db_even.mem_bank[255]);
$fdisplay(file, "0x2000,0x%h_0x%h", db_odd.mem_bank[256],db_even.mem_bank[256]);
$fdisplay(file, "0x2020,0x%h_0x%h", db_odd.mem_bank[257],db_even.mem_bank[257]);
$fdisplay(file, "0x2040,0x%h_0x%h", db_odd.mem_bank[258],db_even.mem_bank[258]);
$fdisplay(file, "0x2060,0x%h_0x%h", db_odd.mem_bank[259],db_even.mem_bank[259]);
$fdisplay(file, "0x2080,0x%h_0x%h", db_odd.mem_bank[260],db_even.mem_bank[260]);
$fdisplay(file, "0x20A0,0x%h_0x%h", db_odd.mem_bank[261],db_even.mem_bank[261]);
$fdisplay(file, "0x20C0,0x%h_0x%h", db_odd.mem_bank[262],db_even.mem_bank[262]);
$fdisplay(file, "0x20E0,0x%h_0x%h", db_odd.mem_bank[263],db_even.mem_bank[263]);
$fdisplay(file, "0x2100,0x%h_0x%h", db_odd.mem_bank[264],db_even.mem_bank[264]);
$fdisplay(file, "0x2120,0x%h_0x%h", db_odd.mem_bank[265],db_even.mem_bank[265]);
$fdisplay(file, "0x2140,0x%h_0x%h", db_odd.mem_bank[266],db_even.mem_bank[266]);
$fdisplay(file, "0x2160,0x%h_0x%h", db_odd.mem_bank[267],db_even.mem_bank[267]);
$fdisplay(file, "0x2180,0x%h_0x%h", db_odd.mem_bank[268],db_even.mem_bank[268]);
$fdisplay(file, "0x21A0,0x%h_0x%h", db_odd.mem_bank[269],db_even.mem_bank[269]);
$fdisplay(file, "0x21C0,0x%h_0x%h", db_odd.mem_bank[270],db_even.mem_bank[270]);
$fdisplay(file, "0x21E0,0x%h_0x%h", db_odd.mem_bank[271],db_even.mem_bank[271]);
$fdisplay(file, "0x2200,0x%h_0x%h", db_odd.mem_bank[272],db_even.mem_bank[272]);
$fdisplay(file, "0x2220,0x%h_0x%h", db_odd.mem_bank[273],db_even.mem_bank[273]);
$fdisplay(file, "0x2240,0x%h_0x%h", db_odd.mem_bank[274],db_even.mem_bank[274]);
$fdisplay(file, "0x2260,0x%h_0x%h", db_odd.mem_bank[275],db_even.mem_bank[275]);
$fdisplay(file, "0x2280,0x%h_0x%h", db_odd.mem_bank[276],db_even.mem_bank[276]);
$fdisplay(file, "0x22A0,0x%h_0x%h", db_odd.mem_bank[277],db_even.mem_bank[277]);
$fdisplay(file, "0x22C0,0x%h_0x%h", db_odd.mem_bank[278],db_even.mem_bank[278]);
$fdisplay(file, "0x22E0,0x%h_0x%h", db_odd.mem_bank[279],db_even.mem_bank[279]);
$fdisplay(file, "0x2300,0x%h_0x%h", db_odd.mem_bank[280],db_even.mem_bank[280]);
$fdisplay(file, "0x2320,0x%h_0x%h", db_odd.mem_bank[281],db_even.mem_bank[281]);
$fdisplay(file, "0x2340,0x%h_0x%h", db_odd.mem_bank[282],db_even.mem_bank[282]);
$fdisplay(file, "0x2360,0x%h_0x%h", db_odd.mem_bank[283],db_even.mem_bank[283]);
$fdisplay(file, "0x2380,0x%h_0x%h", db_odd.mem_bank[284],db_even.mem_bank[284]);
$fdisplay(file, "0x23A0,0x%h_0x%h", db_odd.mem_bank[285],db_even.mem_bank[285]);
$fdisplay(file, "0x23C0,0x%h_0x%h", db_odd.mem_bank[286],db_even.mem_bank[286]);
$fdisplay(file, "0x23E0,0x%h_0x%h", db_odd.mem_bank[287],db_even.mem_bank[287]);
$fdisplay(file, "0x2400,0x%h_0x%h", db_odd.mem_bank[288],db_even.mem_bank[288]);
$fdisplay(file, "0x2420,0x%h_0x%h", db_odd.mem_bank[289],db_even.mem_bank[289]);
$fdisplay(file, "0x2440,0x%h_0x%h", db_odd.mem_bank[290],db_even.mem_bank[290]);
$fdisplay(file, "0x2460,0x%h_0x%h", db_odd.mem_bank[291],db_even.mem_bank[291]);
$fdisplay(file, "0x2480,0x%h_0x%h", db_odd.mem_bank[292],db_even.mem_bank[292]);
$fdisplay(file, "0x24A0,0x%h_0x%h", db_odd.mem_bank[293],db_even.mem_bank[293]);
$fdisplay(file, "0x24C0,0x%h_0x%h", db_odd.mem_bank[294],db_even.mem_bank[294]);
$fdisplay(file, "0x24E0,0x%h_0x%h", db_odd.mem_bank[295],db_even.mem_bank[295]);
$fdisplay(file, "0x2500,0x%h_0x%h", db_odd.mem_bank[296],db_even.mem_bank[296]);
$fdisplay(file, "0x2520,0x%h_0x%h", db_odd.mem_bank[297],db_even.mem_bank[297]);
$fdisplay(file, "0x2540,0x%h_0x%h", db_odd.mem_bank[298],db_even.mem_bank[298]);
$fdisplay(file, "0x2560,0x%h_0x%h", db_odd.mem_bank[299],db_even.mem_bank[299]);
$fdisplay(file, "0x2580,0x%h_0x%h", db_odd.mem_bank[300],db_even.mem_bank[300]);
$fdisplay(file, "0x25A0,0x%h_0x%h", db_odd.mem_bank[301],db_even.mem_bank[301]);
$fdisplay(file, "0x25C0,0x%h_0x%h", db_odd.mem_bank[302],db_even.mem_bank[302]);
$fdisplay(file, "0x25E0,0x%h_0x%h", db_odd.mem_bank[303],db_even.mem_bank[303]);
$fdisplay(file, "0x2600,0x%h_0x%h", db_odd.mem_bank[304],db_even.mem_bank[304]);
$fdisplay(file, "0x2620,0x%h_0x%h", db_odd.mem_bank[305],db_even.mem_bank[305]);
$fdisplay(file, "0x2640,0x%h_0x%h", db_odd.mem_bank[306],db_even.mem_bank[306]);
$fdisplay(file, "0x2660,0x%h_0x%h", db_odd.mem_bank[307],db_even.mem_bank[307]);
$fdisplay(file, "0x2680,0x%h_0x%h", db_odd.mem_bank[308],db_even.mem_bank[308]);
$fdisplay(file, "0x26A0,0x%h_0x%h", db_odd.mem_bank[309],db_even.mem_bank[309]);
$fdisplay(file, "0x26C0,0x%h_0x%h", db_odd.mem_bank[310],db_even.mem_bank[310]);
$fdisplay(file, "0x26E0,0x%h_0x%h", db_odd.mem_bank[311],db_even.mem_bank[311]);
$fdisplay(file, "0x2700,0x%h_0x%h", db_odd.mem_bank[312],db_even.mem_bank[312]);
$fdisplay(file, "0x2720,0x%h_0x%h", db_odd.mem_bank[313],db_even.mem_bank[313]);
$fdisplay(file, "0x2740,0x%h_0x%h", db_odd.mem_bank[314],db_even.mem_bank[314]);
$fdisplay(file, "0x2760,0x%h_0x%h", db_odd.mem_bank[315],db_even.mem_bank[315]);
$fdisplay(file, "0x2780,0x%h_0x%h", db_odd.mem_bank[316],db_even.mem_bank[316]);
$fdisplay(file, "0x27A0,0x%h_0x%h", db_odd.mem_bank[317],db_even.mem_bank[317]);
$fdisplay(file, "0x27C0,0x%h_0x%h", db_odd.mem_bank[318],db_even.mem_bank[318]);
$fdisplay(file, "0x27E0,0x%h_0x%h", db_odd.mem_bank[319],db_even.mem_bank[319]);
$fdisplay(file, "0x2800,0x%h_0x%h", db_odd.mem_bank[320],db_even.mem_bank[320]);
$fdisplay(file, "0x2820,0x%h_0x%h", db_odd.mem_bank[321],db_even.mem_bank[321]);
$fdisplay(file, "0x2840,0x%h_0x%h", db_odd.mem_bank[322],db_even.mem_bank[322]);
$fdisplay(file, "0x2860,0x%h_0x%h", db_odd.mem_bank[323],db_even.mem_bank[323]);
$fdisplay(file, "0x2880,0x%h_0x%h", db_odd.mem_bank[324],db_even.mem_bank[324]);
$fdisplay(file, "0x28A0,0x%h_0x%h", db_odd.mem_bank[325],db_even.mem_bank[325]);
$fdisplay(file, "0x28C0,0x%h_0x%h", db_odd.mem_bank[326],db_even.mem_bank[326]);
$fdisplay(file, "0x28E0,0x%h_0x%h", db_odd.mem_bank[327],db_even.mem_bank[327]);
$fdisplay(file, "0x2900,0x%h_0x%h", db_odd.mem_bank[328],db_even.mem_bank[328]);
$fdisplay(file, "0x2920,0x%h_0x%h", db_odd.mem_bank[329],db_even.mem_bank[329]);
$fdisplay(file, "0x2940,0x%h_0x%h", db_odd.mem_bank[330],db_even.mem_bank[330]);
$fdisplay(file, "0x2960,0x%h_0x%h", db_odd.mem_bank[331],db_even.mem_bank[331]);
$fdisplay(file, "0x2980,0x%h_0x%h", db_odd.mem_bank[332],db_even.mem_bank[332]);
$fdisplay(file, "0x29A0,0x%h_0x%h", db_odd.mem_bank[333],db_even.mem_bank[333]);
$fdisplay(file, "0x29C0,0x%h_0x%h", db_odd.mem_bank[334],db_even.mem_bank[334]);
$fdisplay(file, "0x29E0,0x%h_0x%h", db_odd.mem_bank[335],db_even.mem_bank[335]);
$fdisplay(file, "0x2A00,0x%h_0x%h", db_odd.mem_bank[336],db_even.mem_bank[336]);
$fdisplay(file, "0x2A20,0x%h_0x%h", db_odd.mem_bank[337],db_even.mem_bank[337]);
$fdisplay(file, "0x2A40,0x%h_0x%h", db_odd.mem_bank[338],db_even.mem_bank[338]);
$fdisplay(file, "0x2A60,0x%h_0x%h", db_odd.mem_bank[339],db_even.mem_bank[339]);
$fdisplay(file, "0x2A80,0x%h_0x%h", db_odd.mem_bank[340],db_even.mem_bank[340]);
$fdisplay(file, "0x2AA0,0x%h_0x%h", db_odd.mem_bank[341],db_even.mem_bank[341]);
$fdisplay(file, "0x2AC0,0x%h_0x%h", db_odd.mem_bank[342],db_even.mem_bank[342]);
$fdisplay(file, "0x2AE0,0x%h_0x%h", db_odd.mem_bank[343],db_even.mem_bank[343]);
$fdisplay(file, "0x2B00,0x%h_0x%h", db_odd.mem_bank[344],db_even.mem_bank[344]);
$fdisplay(file, "0x2B20,0x%h_0x%h", db_odd.mem_bank[345],db_even.mem_bank[345]);
$fdisplay(file, "0x2B40,0x%h_0x%h", db_odd.mem_bank[346],db_even.mem_bank[346]);
$fdisplay(file, "0x2B60,0x%h_0x%h", db_odd.mem_bank[347],db_even.mem_bank[347]);
$fdisplay(file, "0x2B80,0x%h_0x%h", db_odd.mem_bank[348],db_even.mem_bank[348]);
$fdisplay(file, "0x2BA0,0x%h_0x%h", db_odd.mem_bank[349],db_even.mem_bank[349]);
$fdisplay(file, "0x2BC0,0x%h_0x%h", db_odd.mem_bank[350],db_even.mem_bank[350]);
$fdisplay(file, "0x2BE0,0x%h_0x%h", db_odd.mem_bank[351],db_even.mem_bank[351]);
$fdisplay(file, "0x2C00,0x%h_0x%h", db_odd.mem_bank[352],db_even.mem_bank[352]);
$fdisplay(file, "0x2C20,0x%h_0x%h", db_odd.mem_bank[353],db_even.mem_bank[353]);
$fdisplay(file, "0x2C40,0x%h_0x%h", db_odd.mem_bank[354],db_even.mem_bank[354]);
$fdisplay(file, "0x2C60,0x%h_0x%h", db_odd.mem_bank[355],db_even.mem_bank[355]);
$fdisplay(file, "0x2C80,0x%h_0x%h", db_odd.mem_bank[356],db_even.mem_bank[356]);
$fdisplay(file, "0x2CA0,0x%h_0x%h", db_odd.mem_bank[357],db_even.mem_bank[357]);
$fdisplay(file, "0x2CC0,0x%h_0x%h", db_odd.mem_bank[358],db_even.mem_bank[358]);
$fdisplay(file, "0x2CE0,0x%h_0x%h", db_odd.mem_bank[359],db_even.mem_bank[359]);
$fdisplay(file, "0x2D00,0x%h_0x%h", db_odd.mem_bank[360],db_even.mem_bank[360]);
$fdisplay(file, "0x2D20,0x%h_0x%h", db_odd.mem_bank[361],db_even.mem_bank[361]);
$fdisplay(file, "0x2D40,0x%h_0x%h", db_odd.mem_bank[362],db_even.mem_bank[362]);
$fdisplay(file, "0x2D60,0x%h_0x%h", db_odd.mem_bank[363],db_even.mem_bank[363]);
$fdisplay(file, "0x2D80,0x%h_0x%h", db_odd.mem_bank[364],db_even.mem_bank[364]);
$fdisplay(file, "0x2DA0,0x%h_0x%h", db_odd.mem_bank[365],db_even.mem_bank[365]);
$fdisplay(file, "0x2DC0,0x%h_0x%h", db_odd.mem_bank[366],db_even.mem_bank[366]);
$fdisplay(file, "0x2DE0,0x%h_0x%h", db_odd.mem_bank[367],db_even.mem_bank[367]);
$fdisplay(file, "0x2E00,0x%h_0x%h", db_odd.mem_bank[368],db_even.mem_bank[368]);
$fdisplay(file, "0x2E20,0x%h_0x%h", db_odd.mem_bank[369],db_even.mem_bank[369]);
$fdisplay(file, "0x2E40,0x%h_0x%h", db_odd.mem_bank[370],db_even.mem_bank[370]);
$fdisplay(file, "0x2E60,0x%h_0x%h", db_odd.mem_bank[371],db_even.mem_bank[371]);
$fdisplay(file, "0x2E80,0x%h_0x%h", db_odd.mem_bank[372],db_even.mem_bank[372]);
$fdisplay(file, "0x2EA0,0x%h_0x%h", db_odd.mem_bank[373],db_even.mem_bank[373]);
$fdisplay(file, "0x2EC0,0x%h_0x%h", db_odd.mem_bank[374],db_even.mem_bank[374]);
$fdisplay(file, "0x2EE0,0x%h_0x%h", db_odd.mem_bank[375],db_even.mem_bank[375]);
$fdisplay(file, "0x2F00,0x%h_0x%h", db_odd.mem_bank[376],db_even.mem_bank[376]);
$fdisplay(file, "0x2F20,0x%h_0x%h", db_odd.mem_bank[377],db_even.mem_bank[377]);
$fdisplay(file, "0x2F40,0x%h_0x%h", db_odd.mem_bank[378],db_even.mem_bank[378]);
$fdisplay(file, "0x2F60,0x%h_0x%h", db_odd.mem_bank[379],db_even.mem_bank[379]);
$fdisplay(file, "0x2F80,0x%h_0x%h", db_odd.mem_bank[380],db_even.mem_bank[380]);
$fdisplay(file, "0x2FA0,0x%h_0x%h", db_odd.mem_bank[381],db_even.mem_bank[381]);
$fdisplay(file, "0x2FC0,0x%h_0x%h", db_odd.mem_bank[382],db_even.mem_bank[382]);
$fdisplay(file, "0x2FE0,0x%h_0x%h", db_odd.mem_bank[383],db_even.mem_bank[383]);
$fdisplay(file, "0x3000,0x%h_0x%h", db_odd.mem_bank[384],db_even.mem_bank[384]);
$fdisplay(file, "0x3020,0x%h_0x%h", db_odd.mem_bank[385],db_even.mem_bank[385]);
$fdisplay(file, "0x3040,0x%h_0x%h", db_odd.mem_bank[386],db_even.mem_bank[386]);
$fdisplay(file, "0x3060,0x%h_0x%h", db_odd.mem_bank[387],db_even.mem_bank[387]);
$fdisplay(file, "0x3080,0x%h_0x%h", db_odd.mem_bank[388],db_even.mem_bank[388]);
$fdisplay(file, "0x30A0,0x%h_0x%h", db_odd.mem_bank[389],db_even.mem_bank[389]);
$fdisplay(file, "0x30C0,0x%h_0x%h", db_odd.mem_bank[390],db_even.mem_bank[390]);
$fdisplay(file, "0x30E0,0x%h_0x%h", db_odd.mem_bank[391],db_even.mem_bank[391]);
$fdisplay(file, "0x3100,0x%h_0x%h", db_odd.mem_bank[392],db_even.mem_bank[392]);
$fdisplay(file, "0x3120,0x%h_0x%h", db_odd.mem_bank[393],db_even.mem_bank[393]);
$fdisplay(file, "0x3140,0x%h_0x%h", db_odd.mem_bank[394],db_even.mem_bank[394]);
$fdisplay(file, "0x3160,0x%h_0x%h", db_odd.mem_bank[395],db_even.mem_bank[395]);
$fdisplay(file, "0x3180,0x%h_0x%h", db_odd.mem_bank[396],db_even.mem_bank[396]);
$fdisplay(file, "0x31A0,0x%h_0x%h", db_odd.mem_bank[397],db_even.mem_bank[397]);
$fdisplay(file, "0x31C0,0x%h_0x%h", db_odd.mem_bank[398],db_even.mem_bank[398]);
$fdisplay(file, "0x31E0,0x%h_0x%h", db_odd.mem_bank[399],db_even.mem_bank[399]);
$fdisplay(file, "0x3200,0x%h_0x%h", db_odd.mem_bank[400],db_even.mem_bank[400]);
$fdisplay(file, "0x3220,0x%h_0x%h", db_odd.mem_bank[401],db_even.mem_bank[401]);
$fdisplay(file, "0x3240,0x%h_0x%h", db_odd.mem_bank[402],db_even.mem_bank[402]);
$fdisplay(file, "0x3260,0x%h_0x%h", db_odd.mem_bank[403],db_even.mem_bank[403]);
$fdisplay(file, "0x3280,0x%h_0x%h", db_odd.mem_bank[404],db_even.mem_bank[404]);
$fdisplay(file, "0x32A0,0x%h_0x%h", db_odd.mem_bank[405],db_even.mem_bank[405]);
$fdisplay(file, "0x32C0,0x%h_0x%h", db_odd.mem_bank[406],db_even.mem_bank[406]);
$fdisplay(file, "0x32E0,0x%h_0x%h", db_odd.mem_bank[407],db_even.mem_bank[407]);
$fdisplay(file, "0x3300,0x%h_0x%h", db_odd.mem_bank[408],db_even.mem_bank[408]);
$fdisplay(file, "0x3320,0x%h_0x%h", db_odd.mem_bank[409],db_even.mem_bank[409]);
$fdisplay(file, "0x3340,0x%h_0x%h", db_odd.mem_bank[410],db_even.mem_bank[410]);
$fdisplay(file, "0x3360,0x%h_0x%h", db_odd.mem_bank[411],db_even.mem_bank[411]);
$fdisplay(file, "0x3380,0x%h_0x%h", db_odd.mem_bank[412],db_even.mem_bank[412]);
$fdisplay(file, "0x33A0,0x%h_0x%h", db_odd.mem_bank[413],db_even.mem_bank[413]);
$fdisplay(file, "0x33C0,0x%h_0x%h", db_odd.mem_bank[414],db_even.mem_bank[414]);
$fdisplay(file, "0x33E0,0x%h_0x%h", db_odd.mem_bank[415],db_even.mem_bank[415]);
$fdisplay(file, "0x3400,0x%h_0x%h", db_odd.mem_bank[416],db_even.mem_bank[416]);
$fdisplay(file, "0x3420,0x%h_0x%h", db_odd.mem_bank[417],db_even.mem_bank[417]);
$fdisplay(file, "0x3440,0x%h_0x%h", db_odd.mem_bank[418],db_even.mem_bank[418]);
$fdisplay(file, "0x3460,0x%h_0x%h", db_odd.mem_bank[419],db_even.mem_bank[419]);
$fdisplay(file, "0x3480,0x%h_0x%h", db_odd.mem_bank[420],db_even.mem_bank[420]);
$fdisplay(file, "0x34A0,0x%h_0x%h", db_odd.mem_bank[421],db_even.mem_bank[421]);
$fdisplay(file, "0x34C0,0x%h_0x%h", db_odd.mem_bank[422],db_even.mem_bank[422]);
$fdisplay(file, "0x34E0,0x%h_0x%h", db_odd.mem_bank[423],db_even.mem_bank[423]);
$fdisplay(file, "0x3500,0x%h_0x%h", db_odd.mem_bank[424],db_even.mem_bank[424]);
$fdisplay(file, "0x3520,0x%h_0x%h", db_odd.mem_bank[425],db_even.mem_bank[425]);
$fdisplay(file, "0x3540,0x%h_0x%h", db_odd.mem_bank[426],db_even.mem_bank[426]);
$fdisplay(file, "0x3560,0x%h_0x%h", db_odd.mem_bank[427],db_even.mem_bank[427]);
$fdisplay(file, "0x3580,0x%h_0x%h", db_odd.mem_bank[428],db_even.mem_bank[428]);
$fdisplay(file, "0x35A0,0x%h_0x%h", db_odd.mem_bank[429],db_even.mem_bank[429]);
$fdisplay(file, "0x35C0,0x%h_0x%h", db_odd.mem_bank[430],db_even.mem_bank[430]);
$fdisplay(file, "0x35E0,0x%h_0x%h", db_odd.mem_bank[431],db_even.mem_bank[431]);
$fdisplay(file, "0x3600,0x%h_0x%h", db_odd.mem_bank[432],db_even.mem_bank[432]);
$fdisplay(file, "0x3620,0x%h_0x%h", db_odd.mem_bank[433],db_even.mem_bank[433]);
$fdisplay(file, "0x3640,0x%h_0x%h", db_odd.mem_bank[434],db_even.mem_bank[434]);
$fdisplay(file, "0x3660,0x%h_0x%h", db_odd.mem_bank[435],db_even.mem_bank[435]);
$fdisplay(file, "0x3680,0x%h_0x%h", db_odd.mem_bank[436],db_even.mem_bank[436]);
$fdisplay(file, "0x36A0,0x%h_0x%h", db_odd.mem_bank[437],db_even.mem_bank[437]);
$fdisplay(file, "0x36C0,0x%h_0x%h", db_odd.mem_bank[438],db_even.mem_bank[438]);
$fdisplay(file, "0x36E0,0x%h_0x%h", db_odd.mem_bank[439],db_even.mem_bank[439]);
$fdisplay(file, "0x3700,0x%h_0x%h", db_odd.mem_bank[440],db_even.mem_bank[440]);
$fdisplay(file, "0x3720,0x%h_0x%h", db_odd.mem_bank[441],db_even.mem_bank[441]);
$fdisplay(file, "0x3740,0x%h_0x%h", db_odd.mem_bank[442],db_even.mem_bank[442]);
$fdisplay(file, "0x3760,0x%h_0x%h", db_odd.mem_bank[443],db_even.mem_bank[443]);
$fdisplay(file, "0x3780,0x%h_0x%h", db_odd.mem_bank[444],db_even.mem_bank[444]);
$fdisplay(file, "0x37A0,0x%h_0x%h", db_odd.mem_bank[445],db_even.mem_bank[445]);
$fdisplay(file, "0x37C0,0x%h_0x%h", db_odd.mem_bank[446],db_even.mem_bank[446]);
$fdisplay(file, "0x37E0,0x%h_0x%h", db_odd.mem_bank[447],db_even.mem_bank[447]);
$fdisplay(file, "0x3800,0x%h_0x%h", db_odd.mem_bank[448],db_even.mem_bank[448]);
$fdisplay(file, "0x3820,0x%h_0x%h", db_odd.mem_bank[449],db_even.mem_bank[449]);
$fdisplay(file, "0x3840,0x%h_0x%h", db_odd.mem_bank[450],db_even.mem_bank[450]);
$fdisplay(file, "0x3860,0x%h_0x%h", db_odd.mem_bank[451],db_even.mem_bank[451]);
$fdisplay(file, "0x3880,0x%h_0x%h", db_odd.mem_bank[452],db_even.mem_bank[452]);
$fdisplay(file, "0x38A0,0x%h_0x%h", db_odd.mem_bank[453],db_even.mem_bank[453]);
$fdisplay(file, "0x38C0,0x%h_0x%h", db_odd.mem_bank[454],db_even.mem_bank[454]);
$fdisplay(file, "0x38E0,0x%h_0x%h", db_odd.mem_bank[455],db_even.mem_bank[455]);
$fdisplay(file, "0x3900,0x%h_0x%h", db_odd.mem_bank[456],db_even.mem_bank[456]);
$fdisplay(file, "0x3920,0x%h_0x%h", db_odd.mem_bank[457],db_even.mem_bank[457]);
$fdisplay(file, "0x3940,0x%h_0x%h", db_odd.mem_bank[458],db_even.mem_bank[458]);
$fdisplay(file, "0x3960,0x%h_0x%h", db_odd.mem_bank[459],db_even.mem_bank[459]);
$fdisplay(file, "0x3980,0x%h_0x%h", db_odd.mem_bank[460],db_even.mem_bank[460]);
$fdisplay(file, "0x39A0,0x%h_0x%h", db_odd.mem_bank[461],db_even.mem_bank[461]);
$fdisplay(file, "0x39C0,0x%h_0x%h", db_odd.mem_bank[462],db_even.mem_bank[462]);
$fdisplay(file, "0x39E0,0x%h_0x%h", db_odd.mem_bank[463],db_even.mem_bank[463]);
$fdisplay(file, "0x3A00,0x%h_0x%h", db_odd.mem_bank[464],db_even.mem_bank[464]);
$fdisplay(file, "0x3A20,0x%h_0x%h", db_odd.mem_bank[465],db_even.mem_bank[465]);
$fdisplay(file, "0x3A40,0x%h_0x%h", db_odd.mem_bank[466],db_even.mem_bank[466]);
$fdisplay(file, "0x3A60,0x%h_0x%h", db_odd.mem_bank[467],db_even.mem_bank[467]);
$fdisplay(file, "0x3A80,0x%h_0x%h", db_odd.mem_bank[468],db_even.mem_bank[468]);
$fdisplay(file, "0x3AA0,0x%h_0x%h", db_odd.mem_bank[469],db_even.mem_bank[469]);
$fdisplay(file, "0x3AC0,0x%h_0x%h", db_odd.mem_bank[470],db_even.mem_bank[470]);
$fdisplay(file, "0x3AE0,0x%h_0x%h", db_odd.mem_bank[471],db_even.mem_bank[471]);
$fdisplay(file, "0x3B00,0x%h_0x%h", db_odd.mem_bank[472],db_even.mem_bank[472]);
$fdisplay(file, "0x3B20,0x%h_0x%h", db_odd.mem_bank[473],db_even.mem_bank[473]);
$fdisplay(file, "0x3B40,0x%h_0x%h", db_odd.mem_bank[474],db_even.mem_bank[474]);
$fdisplay(file, "0x3B60,0x%h_0x%h", db_odd.mem_bank[475],db_even.mem_bank[475]);
$fdisplay(file, "0x3B80,0x%h_0x%h", db_odd.mem_bank[476],db_even.mem_bank[476]);
$fdisplay(file, "0x3BA0,0x%h_0x%h", db_odd.mem_bank[477],db_even.mem_bank[477]);
$fdisplay(file, "0x3BC0,0x%h_0x%h", db_odd.mem_bank[478],db_even.mem_bank[478]);
$fdisplay(file, "0x3BE0,0x%h_0x%h", db_odd.mem_bank[479],db_even.mem_bank[479]);
$fdisplay(file, "0x3C00,0x%h_0x%h", db_odd.mem_bank[480],db_even.mem_bank[480]);
$fdisplay(file, "0x3C20,0x%h_0x%h", db_odd.mem_bank[481],db_even.mem_bank[481]);
$fdisplay(file, "0x3C40,0x%h_0x%h", db_odd.mem_bank[482],db_even.mem_bank[482]);
$fdisplay(file, "0x3C60,0x%h_0x%h", db_odd.mem_bank[483],db_even.mem_bank[483]);
$fdisplay(file, "0x3C80,0x%h_0x%h", db_odd.mem_bank[484],db_even.mem_bank[484]);
$fdisplay(file, "0x3CA0,0x%h_0x%h", db_odd.mem_bank[485],db_even.mem_bank[485]);
$fdisplay(file, "0x3CC0,0x%h_0x%h", db_odd.mem_bank[486],db_even.mem_bank[486]);
$fdisplay(file, "0x3CE0,0x%h_0x%h", db_odd.mem_bank[487],db_even.mem_bank[487]);
$fdisplay(file, "0x3D00,0x%h_0x%h", db_odd.mem_bank[488],db_even.mem_bank[488]);
$fdisplay(file, "0x3D20,0x%h_0x%h", db_odd.mem_bank[489],db_even.mem_bank[489]);
$fdisplay(file, "0x3D40,0x%h_0x%h", db_odd.mem_bank[490],db_even.mem_bank[490]);
$fdisplay(file, "0x3D60,0x%h_0x%h", db_odd.mem_bank[491],db_even.mem_bank[491]);
$fdisplay(file, "0x3D80,0x%h_0x%h", db_odd.mem_bank[492],db_even.mem_bank[492]);
$fdisplay(file, "0x3DA0,0x%h_0x%h", db_odd.mem_bank[493],db_even.mem_bank[493]);
$fdisplay(file, "0x3DC0,0x%h_0x%h", db_odd.mem_bank[494],db_even.mem_bank[494]);
$fdisplay(file, "0x3DE0,0x%h_0x%h", db_odd.mem_bank[495],db_even.mem_bank[495]);
$fdisplay(file, "0x3E00,0x%h_0x%h", db_odd.mem_bank[496],db_even.mem_bank[496]);
$fdisplay(file, "0x3E20,0x%h_0x%h", db_odd.mem_bank[497],db_even.mem_bank[497]);
$fdisplay(file, "0x3E40,0x%h_0x%h", db_odd.mem_bank[498],db_even.mem_bank[498]);
$fdisplay(file, "0x3E60,0x%h_0x%h", db_odd.mem_bank[499],db_even.mem_bank[499]);
$fdisplay(file, "0x3E80,0x%h_0x%h", db_odd.mem_bank[500],db_even.mem_bank[500]);
$fdisplay(file, "0x3EA0,0x%h_0x%h", db_odd.mem_bank[501],db_even.mem_bank[501]);
$fdisplay(file, "0x3EC0,0x%h_0x%h", db_odd.mem_bank[502],db_even.mem_bank[502]);
$fdisplay(file, "0x3EE0,0x%h_0x%h", db_odd.mem_bank[503],db_even.mem_bank[503]);
$fdisplay(file, "0x3F00,0x%h_0x%h", db_odd.mem_bank[504],db_even.mem_bank[504]);
$fdisplay(file, "0x3F20,0x%h_0x%h", db_odd.mem_bank[505],db_even.mem_bank[505]);
$fdisplay(file, "0x3F40,0x%h_0x%h", db_odd.mem_bank[506],db_even.mem_bank[506]);
$fdisplay(file, "0x3F60,0x%h_0x%h", db_odd.mem_bank[507],db_even.mem_bank[507]);
$fdisplay(file, "0x3F80,0x%h_0x%h", db_odd.mem_bank[508],db_even.mem_bank[508]);
$fdisplay(file, "0x3FA0,0x%h_0x%h", db_odd.mem_bank[509],db_even.mem_bank[509]);
$fdisplay(file, "0x3FC0,0x%h_0x%h", db_odd.mem_bank[510],db_even.mem_bank[510]);
$fdisplay(file, "0x3FE0,0x%h_0x%h", db_odd.mem_bank[511],db_even.mem_bank[511]);
$fdisplay(file, "0x4000,0x%h_0x%h", db_odd.mem_bank[512],db_even.mem_bank[512]);
$fdisplay(file, "0x4020,0x%h_0x%h", db_odd.mem_bank[513],db_even.mem_bank[513]);
$fdisplay(file, "0x4040,0x%h_0x%h", db_odd.mem_bank[514],db_even.mem_bank[514]);
$fdisplay(file, "0x4060,0x%h_0x%h", db_odd.mem_bank[515],db_even.mem_bank[515]);
$fdisplay(file, "0x4080,0x%h_0x%h", db_odd.mem_bank[516],db_even.mem_bank[516]);
$fdisplay(file, "0x40A0,0x%h_0x%h", db_odd.mem_bank[517],db_even.mem_bank[517]);
$fdisplay(file, "0x40C0,0x%h_0x%h", db_odd.mem_bank[518],db_even.mem_bank[518]);
$fdisplay(file, "0x40E0,0x%h_0x%h", db_odd.mem_bank[519],db_even.mem_bank[519]);
$fdisplay(file, "0x4100,0x%h_0x%h", db_odd.mem_bank[520],db_even.mem_bank[520]);
$fdisplay(file, "0x4120,0x%h_0x%h", db_odd.mem_bank[521],db_even.mem_bank[521]);
$fdisplay(file, "0x4140,0x%h_0x%h", db_odd.mem_bank[522],db_even.mem_bank[522]);
$fdisplay(file, "0x4160,0x%h_0x%h", db_odd.mem_bank[523],db_even.mem_bank[523]);
$fdisplay(file, "0x4180,0x%h_0x%h", db_odd.mem_bank[524],db_even.mem_bank[524]);
$fdisplay(file, "0x41A0,0x%h_0x%h", db_odd.mem_bank[525],db_even.mem_bank[525]);
$fdisplay(file, "0x41C0,0x%h_0x%h", db_odd.mem_bank[526],db_even.mem_bank[526]);
$fdisplay(file, "0x41E0,0x%h_0x%h", db_odd.mem_bank[527],db_even.mem_bank[527]);
$fdisplay(file, "0x4200,0x%h_0x%h", db_odd.mem_bank[528],db_even.mem_bank[528]);
$fdisplay(file, "0x4220,0x%h_0x%h", db_odd.mem_bank[529],db_even.mem_bank[529]);
$fdisplay(file, "0x4240,0x%h_0x%h", db_odd.mem_bank[530],db_even.mem_bank[530]);
$fdisplay(file, "0x4260,0x%h_0x%h", db_odd.mem_bank[531],db_even.mem_bank[531]);
$fdisplay(file, "0x4280,0x%h_0x%h", db_odd.mem_bank[532],db_even.mem_bank[532]);
$fdisplay(file, "0x42A0,0x%h_0x%h", db_odd.mem_bank[533],db_even.mem_bank[533]);
$fdisplay(file, "0x42C0,0x%h_0x%h", db_odd.mem_bank[534],db_even.mem_bank[534]);
$fdisplay(file, "0x42E0,0x%h_0x%h", db_odd.mem_bank[535],db_even.mem_bank[535]);
$fdisplay(file, "0x4300,0x%h_0x%h", db_odd.mem_bank[536],db_even.mem_bank[536]);
$fdisplay(file, "0x4320,0x%h_0x%h", db_odd.mem_bank[537],db_even.mem_bank[537]);
$fdisplay(file, "0x4340,0x%h_0x%h", db_odd.mem_bank[538],db_even.mem_bank[538]);
$fdisplay(file, "0x4360,0x%h_0x%h", db_odd.mem_bank[539],db_even.mem_bank[539]);
$fdisplay(file, "0x4380,0x%h_0x%h", db_odd.mem_bank[540],db_even.mem_bank[540]);
$fdisplay(file, "0x43A0,0x%h_0x%h", db_odd.mem_bank[541],db_even.mem_bank[541]);
$fdisplay(file, "0x43C0,0x%h_0x%h", db_odd.mem_bank[542],db_even.mem_bank[542]);
$fdisplay(file, "0x43E0,0x%h_0x%h", db_odd.mem_bank[543],db_even.mem_bank[543]);
$fdisplay(file, "0x4400,0x%h_0x%h", db_odd.mem_bank[544],db_even.mem_bank[544]);
$fdisplay(file, "0x4420,0x%h_0x%h", db_odd.mem_bank[545],db_even.mem_bank[545]);
$fdisplay(file, "0x4440,0x%h_0x%h", db_odd.mem_bank[546],db_even.mem_bank[546]);
$fdisplay(file, "0x4460,0x%h_0x%h", db_odd.mem_bank[547],db_even.mem_bank[547]);
$fdisplay(file, "0x4480,0x%h_0x%h", db_odd.mem_bank[548],db_even.mem_bank[548]);
$fdisplay(file, "0x44A0,0x%h_0x%h", db_odd.mem_bank[549],db_even.mem_bank[549]);
$fdisplay(file, "0x44C0,0x%h_0x%h", db_odd.mem_bank[550],db_even.mem_bank[550]);
$fdisplay(file, "0x44E0,0x%h_0x%h", db_odd.mem_bank[551],db_even.mem_bank[551]);
$fdisplay(file, "0x4500,0x%h_0x%h", db_odd.mem_bank[552],db_even.mem_bank[552]);
$fdisplay(file, "0x4520,0x%h_0x%h", db_odd.mem_bank[553],db_even.mem_bank[553]);
$fdisplay(file, "0x4540,0x%h_0x%h", db_odd.mem_bank[554],db_even.mem_bank[554]);
$fdisplay(file, "0x4560,0x%h_0x%h", db_odd.mem_bank[555],db_even.mem_bank[555]);
$fdisplay(file, "0x4580,0x%h_0x%h", db_odd.mem_bank[556],db_even.mem_bank[556]);
$fdisplay(file, "0x45A0,0x%h_0x%h", db_odd.mem_bank[557],db_even.mem_bank[557]);
$fdisplay(file, "0x45C0,0x%h_0x%h", db_odd.mem_bank[558],db_even.mem_bank[558]);
$fdisplay(file, "0x45E0,0x%h_0x%h", db_odd.mem_bank[559],db_even.mem_bank[559]);
$fdisplay(file, "0x4600,0x%h_0x%h", db_odd.mem_bank[560],db_even.mem_bank[560]);
$fdisplay(file, "0x4620,0x%h_0x%h", db_odd.mem_bank[561],db_even.mem_bank[561]);
$fdisplay(file, "0x4640,0x%h_0x%h", db_odd.mem_bank[562],db_even.mem_bank[562]);
$fdisplay(file, "0x4660,0x%h_0x%h", db_odd.mem_bank[563],db_even.mem_bank[563]);
$fdisplay(file, "0x4680,0x%h_0x%h", db_odd.mem_bank[564],db_even.mem_bank[564]);
$fdisplay(file, "0x46A0,0x%h_0x%h", db_odd.mem_bank[565],db_even.mem_bank[565]);
$fdisplay(file, "0x46C0,0x%h_0x%h", db_odd.mem_bank[566],db_even.mem_bank[566]);
$fdisplay(file, "0x46E0,0x%h_0x%h", db_odd.mem_bank[567],db_even.mem_bank[567]);
$fdisplay(file, "0x4700,0x%h_0x%h", db_odd.mem_bank[568],db_even.mem_bank[568]);
$fdisplay(file, "0x4720,0x%h_0x%h", db_odd.mem_bank[569],db_even.mem_bank[569]);
$fdisplay(file, "0x4740,0x%h_0x%h", db_odd.mem_bank[570],db_even.mem_bank[570]);
$fdisplay(file, "0x4760,0x%h_0x%h", db_odd.mem_bank[571],db_even.mem_bank[571]);
$fdisplay(file, "0x4780,0x%h_0x%h", db_odd.mem_bank[572],db_even.mem_bank[572]);
$fdisplay(file, "0x47A0,0x%h_0x%h", db_odd.mem_bank[573],db_even.mem_bank[573]);
$fdisplay(file, "0x47C0,0x%h_0x%h", db_odd.mem_bank[574],db_even.mem_bank[574]);
$fdisplay(file, "0x47E0,0x%h_0x%h", db_odd.mem_bank[575],db_even.mem_bank[575]);
$fdisplay(file, "0x4800,0x%h_0x%h", db_odd.mem_bank[576],db_even.mem_bank[576]);
$fdisplay(file, "0x4820,0x%h_0x%h", db_odd.mem_bank[577],db_even.mem_bank[577]);
$fdisplay(file, "0x4840,0x%h_0x%h", db_odd.mem_bank[578],db_even.mem_bank[578]);
$fdisplay(file, "0x4860,0x%h_0x%h", db_odd.mem_bank[579],db_even.mem_bank[579]);
$fdisplay(file, "0x4880,0x%h_0x%h", db_odd.mem_bank[580],db_even.mem_bank[580]);
$fdisplay(file, "0x48A0,0x%h_0x%h", db_odd.mem_bank[581],db_even.mem_bank[581]);
$fdisplay(file, "0x48C0,0x%h_0x%h", db_odd.mem_bank[582],db_even.mem_bank[582]);
$fdisplay(file, "0x48E0,0x%h_0x%h", db_odd.mem_bank[583],db_even.mem_bank[583]);
$fdisplay(file, "0x4900,0x%h_0x%h", db_odd.mem_bank[584],db_even.mem_bank[584]);
$fdisplay(file, "0x4920,0x%h_0x%h", db_odd.mem_bank[585],db_even.mem_bank[585]);
$fdisplay(file, "0x4940,0x%h_0x%h", db_odd.mem_bank[586],db_even.mem_bank[586]);
$fdisplay(file, "0x4960,0x%h_0x%h", db_odd.mem_bank[587],db_even.mem_bank[587]);
$fdisplay(file, "0x4980,0x%h_0x%h", db_odd.mem_bank[588],db_even.mem_bank[588]);
$fdisplay(file, "0x49A0,0x%h_0x%h", db_odd.mem_bank[589],db_even.mem_bank[589]);
$fdisplay(file, "0x49C0,0x%h_0x%h", db_odd.mem_bank[590],db_even.mem_bank[590]);
$fdisplay(file, "0x49E0,0x%h_0x%h", db_odd.mem_bank[591],db_even.mem_bank[591]);
$fdisplay(file, "0x4A00,0x%h_0x%h", db_odd.mem_bank[592],db_even.mem_bank[592]);
$fdisplay(file, "0x4A20,0x%h_0x%h", db_odd.mem_bank[593],db_even.mem_bank[593]);
$fdisplay(file, "0x4A40,0x%h_0x%h", db_odd.mem_bank[594],db_even.mem_bank[594]);
$fdisplay(file, "0x4A60,0x%h_0x%h", db_odd.mem_bank[595],db_even.mem_bank[595]);
$fdisplay(file, "0x4A80,0x%h_0x%h", db_odd.mem_bank[596],db_even.mem_bank[596]);
$fdisplay(file, "0x4AA0,0x%h_0x%h", db_odd.mem_bank[597],db_even.mem_bank[597]);
$fdisplay(file, "0x4AC0,0x%h_0x%h", db_odd.mem_bank[598],db_even.mem_bank[598]);
$fdisplay(file, "0x4AE0,0x%h_0x%h", db_odd.mem_bank[599],db_even.mem_bank[599]);
$fdisplay(file, "0x4B00,0x%h_0x%h", db_odd.mem_bank[600],db_even.mem_bank[600]);
$fdisplay(file, "0x4B20,0x%h_0x%h", db_odd.mem_bank[601],db_even.mem_bank[601]);
$fdisplay(file, "0x4B40,0x%h_0x%h", db_odd.mem_bank[602],db_even.mem_bank[602]);
$fdisplay(file, "0x4B60,0x%h_0x%h", db_odd.mem_bank[603],db_even.mem_bank[603]);
$fdisplay(file, "0x4B80,0x%h_0x%h", db_odd.mem_bank[604],db_even.mem_bank[604]);
$fdisplay(file, "0x4BA0,0x%h_0x%h", db_odd.mem_bank[605],db_even.mem_bank[605]);
$fdisplay(file, "0x4BC0,0x%h_0x%h", db_odd.mem_bank[606],db_even.mem_bank[606]);
$fdisplay(file, "0x4BE0,0x%h_0x%h", db_odd.mem_bank[607],db_even.mem_bank[607]);
$fdisplay(file, "0x4C00,0x%h_0x%h", db_odd.mem_bank[608],db_even.mem_bank[608]);
$fdisplay(file, "0x4C20,0x%h_0x%h", db_odd.mem_bank[609],db_even.mem_bank[609]);
$fdisplay(file, "0x4C40,0x%h_0x%h", db_odd.mem_bank[610],db_even.mem_bank[610]);
$fdisplay(file, "0x4C60,0x%h_0x%h", db_odd.mem_bank[611],db_even.mem_bank[611]);
$fdisplay(file, "0x4C80,0x%h_0x%h", db_odd.mem_bank[612],db_even.mem_bank[612]);
$fdisplay(file, "0x4CA0,0x%h_0x%h", db_odd.mem_bank[613],db_even.mem_bank[613]);
$fdisplay(file, "0x4CC0,0x%h_0x%h", db_odd.mem_bank[614],db_even.mem_bank[614]);
$fdisplay(file, "0x4CE0,0x%h_0x%h", db_odd.mem_bank[615],db_even.mem_bank[615]);
$fdisplay(file, "0x4D00,0x%h_0x%h", db_odd.mem_bank[616],db_even.mem_bank[616]);
$fdisplay(file, "0x4D20,0x%h_0x%h", db_odd.mem_bank[617],db_even.mem_bank[617]);
$fdisplay(file, "0x4D40,0x%h_0x%h", db_odd.mem_bank[618],db_even.mem_bank[618]);
$fdisplay(file, "0x4D60,0x%h_0x%h", db_odd.mem_bank[619],db_even.mem_bank[619]);
$fdisplay(file, "0x4D80,0x%h_0x%h", db_odd.mem_bank[620],db_even.mem_bank[620]);
$fdisplay(file, "0x4DA0,0x%h_0x%h", db_odd.mem_bank[621],db_even.mem_bank[621]);
$fdisplay(file, "0x4DC0,0x%h_0x%h", db_odd.mem_bank[622],db_even.mem_bank[622]);
$fdisplay(file, "0x4DE0,0x%h_0x%h", db_odd.mem_bank[623],db_even.mem_bank[623]);
$fdisplay(file, "0x4E00,0x%h_0x%h", db_odd.mem_bank[624],db_even.mem_bank[624]);
$fdisplay(file, "0x4E20,0x%h_0x%h", db_odd.mem_bank[625],db_even.mem_bank[625]);
$fdisplay(file, "0x4E40,0x%h_0x%h", db_odd.mem_bank[626],db_even.mem_bank[626]);
$fdisplay(file, "0x4E60,0x%h_0x%h", db_odd.mem_bank[627],db_even.mem_bank[627]);
$fdisplay(file, "0x4E80,0x%h_0x%h", db_odd.mem_bank[628],db_even.mem_bank[628]);
$fdisplay(file, "0x4EA0,0x%h_0x%h", db_odd.mem_bank[629],db_even.mem_bank[629]);
$fdisplay(file, "0x4EC0,0x%h_0x%h", db_odd.mem_bank[630],db_even.mem_bank[630]);
$fdisplay(file, "0x4EE0,0x%h_0x%h", db_odd.mem_bank[631],db_even.mem_bank[631]);
$fdisplay(file, "0x4F00,0x%h_0x%h", db_odd.mem_bank[632],db_even.mem_bank[632]);
$fdisplay(file, "0x4F20,0x%h_0x%h", db_odd.mem_bank[633],db_even.mem_bank[633]);
$fdisplay(file, "0x4F40,0x%h_0x%h", db_odd.mem_bank[634],db_even.mem_bank[634]);
$fdisplay(file, "0x4F60,0x%h_0x%h", db_odd.mem_bank[635],db_even.mem_bank[635]);
$fdisplay(file, "0x4F80,0x%h_0x%h", db_odd.mem_bank[636],db_even.mem_bank[636]);
$fdisplay(file, "0x4FA0,0x%h_0x%h", db_odd.mem_bank[637],db_even.mem_bank[637]);
$fdisplay(file, "0x4FC0,0x%h_0x%h", db_odd.mem_bank[638],db_even.mem_bank[638]);
$fdisplay(file, "0x4FE0,0x%h_0x%h", db_odd.mem_bank[639],db_even.mem_bank[639]);
$fdisplay(file, "0x5000,0x%h_0x%h", db_odd.mem_bank[640],db_even.mem_bank[640]);
$fdisplay(file, "0x5020,0x%h_0x%h", db_odd.mem_bank[641],db_even.mem_bank[641]);
$fdisplay(file, "0x5040,0x%h_0x%h", db_odd.mem_bank[642],db_even.mem_bank[642]);
$fdisplay(file, "0x5060,0x%h_0x%h", db_odd.mem_bank[643],db_even.mem_bank[643]);
$fdisplay(file, "0x5080,0x%h_0x%h", db_odd.mem_bank[644],db_even.mem_bank[644]);
$fdisplay(file, "0x50A0,0x%h_0x%h", db_odd.mem_bank[645],db_even.mem_bank[645]);
$fdisplay(file, "0x50C0,0x%h_0x%h", db_odd.mem_bank[646],db_even.mem_bank[646]);
$fdisplay(file, "0x50E0,0x%h_0x%h", db_odd.mem_bank[647],db_even.mem_bank[647]);
$fdisplay(file, "0x5100,0x%h_0x%h", db_odd.mem_bank[648],db_even.mem_bank[648]);
$fdisplay(file, "0x5120,0x%h_0x%h", db_odd.mem_bank[649],db_even.mem_bank[649]);
$fdisplay(file, "0x5140,0x%h_0x%h", db_odd.mem_bank[650],db_even.mem_bank[650]);
$fdisplay(file, "0x5160,0x%h_0x%h", db_odd.mem_bank[651],db_even.mem_bank[651]);
$fdisplay(file, "0x5180,0x%h_0x%h", db_odd.mem_bank[652],db_even.mem_bank[652]);
$fdisplay(file, "0x51A0,0x%h_0x%h", db_odd.mem_bank[653],db_even.mem_bank[653]);
$fdisplay(file, "0x51C0,0x%h_0x%h", db_odd.mem_bank[654],db_even.mem_bank[654]);
$fdisplay(file, "0x51E0,0x%h_0x%h", db_odd.mem_bank[655],db_even.mem_bank[655]);
$fdisplay(file, "0x5200,0x%h_0x%h", db_odd.mem_bank[656],db_even.mem_bank[656]);
$fdisplay(file, "0x5220,0x%h_0x%h", db_odd.mem_bank[657],db_even.mem_bank[657]);
$fdisplay(file, "0x5240,0x%h_0x%h", db_odd.mem_bank[658],db_even.mem_bank[658]);
$fdisplay(file, "0x5260,0x%h_0x%h", db_odd.mem_bank[659],db_even.mem_bank[659]);
$fdisplay(file, "0x5280,0x%h_0x%h", db_odd.mem_bank[660],db_even.mem_bank[660]);
$fdisplay(file, "0x52A0,0x%h_0x%h", db_odd.mem_bank[661],db_even.mem_bank[661]);
$fdisplay(file, "0x52C0,0x%h_0x%h", db_odd.mem_bank[662],db_even.mem_bank[662]);
$fdisplay(file, "0x52E0,0x%h_0x%h", db_odd.mem_bank[663],db_even.mem_bank[663]);
$fdisplay(file, "0x5300,0x%h_0x%h", db_odd.mem_bank[664],db_even.mem_bank[664]);
$fdisplay(file, "0x5320,0x%h_0x%h", db_odd.mem_bank[665],db_even.mem_bank[665]);
$fdisplay(file, "0x5340,0x%h_0x%h", db_odd.mem_bank[666],db_even.mem_bank[666]);
$fdisplay(file, "0x5360,0x%h_0x%h", db_odd.mem_bank[667],db_even.mem_bank[667]);
$fdisplay(file, "0x5380,0x%h_0x%h", db_odd.mem_bank[668],db_even.mem_bank[668]);
$fdisplay(file, "0x53A0,0x%h_0x%h", db_odd.mem_bank[669],db_even.mem_bank[669]);
$fdisplay(file, "0x53C0,0x%h_0x%h", db_odd.mem_bank[670],db_even.mem_bank[670]);
$fdisplay(file, "0x53E0,0x%h_0x%h", db_odd.mem_bank[671],db_even.mem_bank[671]);
$fdisplay(file, "0x5400,0x%h_0x%h", db_odd.mem_bank[672],db_even.mem_bank[672]);
$fdisplay(file, "0x5420,0x%h_0x%h", db_odd.mem_bank[673],db_even.mem_bank[673]);
$fdisplay(file, "0x5440,0x%h_0x%h", db_odd.mem_bank[674],db_even.mem_bank[674]);
$fdisplay(file, "0x5460,0x%h_0x%h", db_odd.mem_bank[675],db_even.mem_bank[675]);
$fdisplay(file, "0x5480,0x%h_0x%h", db_odd.mem_bank[676],db_even.mem_bank[676]);
$fdisplay(file, "0x54A0,0x%h_0x%h", db_odd.mem_bank[677],db_even.mem_bank[677]);
$fdisplay(file, "0x54C0,0x%h_0x%h", db_odd.mem_bank[678],db_even.mem_bank[678]);
$fdisplay(file, "0x54E0,0x%h_0x%h", db_odd.mem_bank[679],db_even.mem_bank[679]);
$fdisplay(file, "0x5500,0x%h_0x%h", db_odd.mem_bank[680],db_even.mem_bank[680]);
$fdisplay(file, "0x5520,0x%h_0x%h", db_odd.mem_bank[681],db_even.mem_bank[681]);
$fdisplay(file, "0x5540,0x%h_0x%h", db_odd.mem_bank[682],db_even.mem_bank[682]);
$fdisplay(file, "0x5560,0x%h_0x%h", db_odd.mem_bank[683],db_even.mem_bank[683]);
$fdisplay(file, "0x5580,0x%h_0x%h", db_odd.mem_bank[684],db_even.mem_bank[684]);
$fdisplay(file, "0x55A0,0x%h_0x%h", db_odd.mem_bank[685],db_even.mem_bank[685]);
$fdisplay(file, "0x55C0,0x%h_0x%h", db_odd.mem_bank[686],db_even.mem_bank[686]);
$fdisplay(file, "0x55E0,0x%h_0x%h", db_odd.mem_bank[687],db_even.mem_bank[687]);
$fdisplay(file, "0x5600,0x%h_0x%h", db_odd.mem_bank[688],db_even.mem_bank[688]);
$fdisplay(file, "0x5620,0x%h_0x%h", db_odd.mem_bank[689],db_even.mem_bank[689]);
$fdisplay(file, "0x5640,0x%h_0x%h", db_odd.mem_bank[690],db_even.mem_bank[690]);
$fdisplay(file, "0x5660,0x%h_0x%h", db_odd.mem_bank[691],db_even.mem_bank[691]);
$fdisplay(file, "0x5680,0x%h_0x%h", db_odd.mem_bank[692],db_even.mem_bank[692]);
$fdisplay(file, "0x56A0,0x%h_0x%h", db_odd.mem_bank[693],db_even.mem_bank[693]);
$fdisplay(file, "0x56C0,0x%h_0x%h", db_odd.mem_bank[694],db_even.mem_bank[694]);
$fdisplay(file, "0x56E0,0x%h_0x%h", db_odd.mem_bank[695],db_even.mem_bank[695]);
$fdisplay(file, "0x5700,0x%h_0x%h", db_odd.mem_bank[696],db_even.mem_bank[696]);
$fdisplay(file, "0x5720,0x%h_0x%h", db_odd.mem_bank[697],db_even.mem_bank[697]);
$fdisplay(file, "0x5740,0x%h_0x%h", db_odd.mem_bank[698],db_even.mem_bank[698]);
$fdisplay(file, "0x5760,0x%h_0x%h", db_odd.mem_bank[699],db_even.mem_bank[699]);
$fdisplay(file, "0x5780,0x%h_0x%h", db_odd.mem_bank[700],db_even.mem_bank[700]);
$fdisplay(file, "0x57A0,0x%h_0x%h", db_odd.mem_bank[701],db_even.mem_bank[701]);
$fdisplay(file, "0x57C0,0x%h_0x%h", db_odd.mem_bank[702],db_even.mem_bank[702]);
$fdisplay(file, "0x57E0,0x%h_0x%h", db_odd.mem_bank[703],db_even.mem_bank[703]);
$fdisplay(file, "0x5800,0x%h_0x%h", db_odd.mem_bank[704],db_even.mem_bank[704]);
$fdisplay(file, "0x5820,0x%h_0x%h", db_odd.mem_bank[705],db_even.mem_bank[705]);
$fdisplay(file, "0x5840,0x%h_0x%h", db_odd.mem_bank[706],db_even.mem_bank[706]);
$fdisplay(file, "0x5860,0x%h_0x%h", db_odd.mem_bank[707],db_even.mem_bank[707]);
$fdisplay(file, "0x5880,0x%h_0x%h", db_odd.mem_bank[708],db_even.mem_bank[708]);
$fdisplay(file, "0x58A0,0x%h_0x%h", db_odd.mem_bank[709],db_even.mem_bank[709]);
$fdisplay(file, "0x58C0,0x%h_0x%h", db_odd.mem_bank[710],db_even.mem_bank[710]);
$fdisplay(file, "0x58E0,0x%h_0x%h", db_odd.mem_bank[711],db_even.mem_bank[711]);
$fdisplay(file, "0x5900,0x%h_0x%h", db_odd.mem_bank[712],db_even.mem_bank[712]);
$fdisplay(file, "0x5920,0x%h_0x%h", db_odd.mem_bank[713],db_even.mem_bank[713]);
$fdisplay(file, "0x5940,0x%h_0x%h", db_odd.mem_bank[714],db_even.mem_bank[714]);
$fdisplay(file, "0x5960,0x%h_0x%h", db_odd.mem_bank[715],db_even.mem_bank[715]);
$fdisplay(file, "0x5980,0x%h_0x%h", db_odd.mem_bank[716],db_even.mem_bank[716]);
$fdisplay(file, "0x59A0,0x%h_0x%h", db_odd.mem_bank[717],db_even.mem_bank[717]);
$fdisplay(file, "0x59C0,0x%h_0x%h", db_odd.mem_bank[718],db_even.mem_bank[718]);
$fdisplay(file, "0x59E0,0x%h_0x%h", db_odd.mem_bank[719],db_even.mem_bank[719]);
$fdisplay(file, "0x5A00,0x%h_0x%h", db_odd.mem_bank[720],db_even.mem_bank[720]);
$fdisplay(file, "0x5A20,0x%h_0x%h", db_odd.mem_bank[721],db_even.mem_bank[721]);
$fdisplay(file, "0x5A40,0x%h_0x%h", db_odd.mem_bank[722],db_even.mem_bank[722]);
$fdisplay(file, "0x5A60,0x%h_0x%h", db_odd.mem_bank[723],db_even.mem_bank[723]);
$fdisplay(file, "0x5A80,0x%h_0x%h", db_odd.mem_bank[724],db_even.mem_bank[724]);
$fdisplay(file, "0x5AA0,0x%h_0x%h", db_odd.mem_bank[725],db_even.mem_bank[725]);
$fdisplay(file, "0x5AC0,0x%h_0x%h", db_odd.mem_bank[726],db_even.mem_bank[726]);
$fdisplay(file, "0x5AE0,0x%h_0x%h", db_odd.mem_bank[727],db_even.mem_bank[727]);
$fdisplay(file, "0x5B00,0x%h_0x%h", db_odd.mem_bank[728],db_even.mem_bank[728]);
$fdisplay(file, "0x5B20,0x%h_0x%h", db_odd.mem_bank[729],db_even.mem_bank[729]);
$fdisplay(file, "0x5B40,0x%h_0x%h", db_odd.mem_bank[730],db_even.mem_bank[730]);
$fdisplay(file, "0x5B60,0x%h_0x%h", db_odd.mem_bank[731],db_even.mem_bank[731]);
$fdisplay(file, "0x5B80,0x%h_0x%h", db_odd.mem_bank[732],db_even.mem_bank[732]);
$fdisplay(file, "0x5BA0,0x%h_0x%h", db_odd.mem_bank[733],db_even.mem_bank[733]);
$fdisplay(file, "0x5BC0,0x%h_0x%h", db_odd.mem_bank[734],db_even.mem_bank[734]);
$fdisplay(file, "0x5BE0,0x%h_0x%h", db_odd.mem_bank[735],db_even.mem_bank[735]);
$fdisplay(file, "0x5C00,0x%h_0x%h", db_odd.mem_bank[736],db_even.mem_bank[736]);
$fdisplay(file, "0x5C20,0x%h_0x%h", db_odd.mem_bank[737],db_even.mem_bank[737]);
$fdisplay(file, "0x5C40,0x%h_0x%h", db_odd.mem_bank[738],db_even.mem_bank[738]);
$fdisplay(file, "0x5C60,0x%h_0x%h", db_odd.mem_bank[739],db_even.mem_bank[739]);
$fdisplay(file, "0x5C80,0x%h_0x%h", db_odd.mem_bank[740],db_even.mem_bank[740]);
$fdisplay(file, "0x5CA0,0x%h_0x%h", db_odd.mem_bank[741],db_even.mem_bank[741]);
$fdisplay(file, "0x5CC0,0x%h_0x%h", db_odd.mem_bank[742],db_even.mem_bank[742]);
$fdisplay(file, "0x5CE0,0x%h_0x%h", db_odd.mem_bank[743],db_even.mem_bank[743]);
$fdisplay(file, "0x5D00,0x%h_0x%h", db_odd.mem_bank[744],db_even.mem_bank[744]);
$fdisplay(file, "0x5D20,0x%h_0x%h", db_odd.mem_bank[745],db_even.mem_bank[745]);
$fdisplay(file, "0x5D40,0x%h_0x%h", db_odd.mem_bank[746],db_even.mem_bank[746]);
$fdisplay(file, "0x5D60,0x%h_0x%h", db_odd.mem_bank[747],db_even.mem_bank[747]);
$fdisplay(file, "0x5D80,0x%h_0x%h", db_odd.mem_bank[748],db_even.mem_bank[748]);
$fdisplay(file, "0x5DA0,0x%h_0x%h", db_odd.mem_bank[749],db_even.mem_bank[749]);
$fdisplay(file, "0x5DC0,0x%h_0x%h", db_odd.mem_bank[750],db_even.mem_bank[750]);
$fdisplay(file, "0x5DE0,0x%h_0x%h", db_odd.mem_bank[751],db_even.mem_bank[751]);
$fdisplay(file, "0x5E00,0x%h_0x%h", db_odd.mem_bank[752],db_even.mem_bank[752]);
$fdisplay(file, "0x5E20,0x%h_0x%h", db_odd.mem_bank[753],db_even.mem_bank[753]);
$fdisplay(file, "0x5E40,0x%h_0x%h", db_odd.mem_bank[754],db_even.mem_bank[754]);
$fdisplay(file, "0x5E60,0x%h_0x%h", db_odd.mem_bank[755],db_even.mem_bank[755]);
$fdisplay(file, "0x5E80,0x%h_0x%h", db_odd.mem_bank[756],db_even.mem_bank[756]);
$fdisplay(file, "0x5EA0,0x%h_0x%h", db_odd.mem_bank[757],db_even.mem_bank[757]);
$fdisplay(file, "0x5EC0,0x%h_0x%h", db_odd.mem_bank[758],db_even.mem_bank[758]);
$fdisplay(file, "0x5EE0,0x%h_0x%h", db_odd.mem_bank[759],db_even.mem_bank[759]);
$fdisplay(file, "0x5F00,0x%h_0x%h", db_odd.mem_bank[760],db_even.mem_bank[760]);
$fdisplay(file, "0x5F20,0x%h_0x%h", db_odd.mem_bank[761],db_even.mem_bank[761]);
$fdisplay(file, "0x5F40,0x%h_0x%h", db_odd.mem_bank[762],db_even.mem_bank[762]);
$fdisplay(file, "0x5F60,0x%h_0x%h", db_odd.mem_bank[763],db_even.mem_bank[763]);
$fdisplay(file, "0x5F80,0x%h_0x%h", db_odd.mem_bank[764],db_even.mem_bank[764]);
$fdisplay(file, "0x5FA0,0x%h_0x%h", db_odd.mem_bank[765],db_even.mem_bank[765]);
$fdisplay(file, "0x5FC0,0x%h_0x%h", db_odd.mem_bank[766],db_even.mem_bank[766]);
$fdisplay(file, "0x5FE0,0x%h_0x%h", db_odd.mem_bank[767],db_even.mem_bank[767]);
$fdisplay(file, "0x6000,0x%h_0x%h", db_odd.mem_bank[768],db_even.mem_bank[768]);
$fdisplay(file, "0x6020,0x%h_0x%h", db_odd.mem_bank[769],db_even.mem_bank[769]);
$fdisplay(file, "0x6040,0x%h_0x%h", db_odd.mem_bank[770],db_even.mem_bank[770]);
$fdisplay(file, "0x6060,0x%h_0x%h", db_odd.mem_bank[771],db_even.mem_bank[771]);
$fdisplay(file, "0x6080,0x%h_0x%h", db_odd.mem_bank[772],db_even.mem_bank[772]);
$fdisplay(file, "0x60A0,0x%h_0x%h", db_odd.mem_bank[773],db_even.mem_bank[773]);
$fdisplay(file, "0x60C0,0x%h_0x%h", db_odd.mem_bank[774],db_even.mem_bank[774]);
$fdisplay(file, "0x60E0,0x%h_0x%h", db_odd.mem_bank[775],db_even.mem_bank[775]);
$fdisplay(file, "0x6100,0x%h_0x%h", db_odd.mem_bank[776],db_even.mem_bank[776]);
$fdisplay(file, "0x6120,0x%h_0x%h", db_odd.mem_bank[777],db_even.mem_bank[777]);
$fdisplay(file, "0x6140,0x%h_0x%h", db_odd.mem_bank[778],db_even.mem_bank[778]);
$fdisplay(file, "0x6160,0x%h_0x%h", db_odd.mem_bank[779],db_even.mem_bank[779]);
$fdisplay(file, "0x6180,0x%h_0x%h", db_odd.mem_bank[780],db_even.mem_bank[780]);
$fdisplay(file, "0x61A0,0x%h_0x%h", db_odd.mem_bank[781],db_even.mem_bank[781]);
$fdisplay(file, "0x61C0,0x%h_0x%h", db_odd.mem_bank[782],db_even.mem_bank[782]);
$fdisplay(file, "0x61E0,0x%h_0x%h", db_odd.mem_bank[783],db_even.mem_bank[783]);
$fdisplay(file, "0x6200,0x%h_0x%h", db_odd.mem_bank[784],db_even.mem_bank[784]);
$fdisplay(file, "0x6220,0x%h_0x%h", db_odd.mem_bank[785],db_even.mem_bank[785]);
$fdisplay(file, "0x6240,0x%h_0x%h", db_odd.mem_bank[786],db_even.mem_bank[786]);
$fdisplay(file, "0x6260,0x%h_0x%h", db_odd.mem_bank[787],db_even.mem_bank[787]);
$fdisplay(file, "0x6280,0x%h_0x%h", db_odd.mem_bank[788],db_even.mem_bank[788]);
$fdisplay(file, "0x62A0,0x%h_0x%h", db_odd.mem_bank[789],db_even.mem_bank[789]);
$fdisplay(file, "0x62C0,0x%h_0x%h", db_odd.mem_bank[790],db_even.mem_bank[790]);
$fdisplay(file, "0x62E0,0x%h_0x%h", db_odd.mem_bank[791],db_even.mem_bank[791]);
$fdisplay(file, "0x6300,0x%h_0x%h", db_odd.mem_bank[792],db_even.mem_bank[792]);
$fdisplay(file, "0x6320,0x%h_0x%h", db_odd.mem_bank[793],db_even.mem_bank[793]);
$fdisplay(file, "0x6340,0x%h_0x%h", db_odd.mem_bank[794],db_even.mem_bank[794]);
$fdisplay(file, "0x6360,0x%h_0x%h", db_odd.mem_bank[795],db_even.mem_bank[795]);
$fdisplay(file, "0x6380,0x%h_0x%h", db_odd.mem_bank[796],db_even.mem_bank[796]);
$fdisplay(file, "0x63A0,0x%h_0x%h", db_odd.mem_bank[797],db_even.mem_bank[797]);
$fdisplay(file, "0x63C0,0x%h_0x%h", db_odd.mem_bank[798],db_even.mem_bank[798]);
$fdisplay(file, "0x63E0,0x%h_0x%h", db_odd.mem_bank[799],db_even.mem_bank[799]);
$fdisplay(file, "0x6400,0x%h_0x%h", db_odd.mem_bank[800],db_even.mem_bank[800]);
$fdisplay(file, "0x6420,0x%h_0x%h", db_odd.mem_bank[801],db_even.mem_bank[801]);
$fdisplay(file, "0x6440,0x%h_0x%h", db_odd.mem_bank[802],db_even.mem_bank[802]);
$fdisplay(file, "0x6460,0x%h_0x%h", db_odd.mem_bank[803],db_even.mem_bank[803]);
$fdisplay(file, "0x6480,0x%h_0x%h", db_odd.mem_bank[804],db_even.mem_bank[804]);
$fdisplay(file, "0x64A0,0x%h_0x%h", db_odd.mem_bank[805],db_even.mem_bank[805]);
$fdisplay(file, "0x64C0,0x%h_0x%h", db_odd.mem_bank[806],db_even.mem_bank[806]);
$fdisplay(file, "0x64E0,0x%h_0x%h", db_odd.mem_bank[807],db_even.mem_bank[807]);
$fdisplay(file, "0x6500,0x%h_0x%h", db_odd.mem_bank[808],db_even.mem_bank[808]);
$fdisplay(file, "0x6520,0x%h_0x%h", db_odd.mem_bank[809],db_even.mem_bank[809]);
$fdisplay(file, "0x6540,0x%h_0x%h", db_odd.mem_bank[810],db_even.mem_bank[810]);
$fdisplay(file, "0x6560,0x%h_0x%h", db_odd.mem_bank[811],db_even.mem_bank[811]);
$fdisplay(file, "0x6580,0x%h_0x%h", db_odd.mem_bank[812],db_even.mem_bank[812]);
$fdisplay(file, "0x65A0,0x%h_0x%h", db_odd.mem_bank[813],db_even.mem_bank[813]);
$fdisplay(file, "0x65C0,0x%h_0x%h", db_odd.mem_bank[814],db_even.mem_bank[814]);
$fdisplay(file, "0x65E0,0x%h_0x%h", db_odd.mem_bank[815],db_even.mem_bank[815]);
$fdisplay(file, "0x6600,0x%h_0x%h", db_odd.mem_bank[816],db_even.mem_bank[816]);
$fdisplay(file, "0x6620,0x%h_0x%h", db_odd.mem_bank[817],db_even.mem_bank[817]);
$fdisplay(file, "0x6640,0x%h_0x%h", db_odd.mem_bank[818],db_even.mem_bank[818]);
$fdisplay(file, "0x6660,0x%h_0x%h", db_odd.mem_bank[819],db_even.mem_bank[819]);
$fdisplay(file, "0x6680,0x%h_0x%h", db_odd.mem_bank[820],db_even.mem_bank[820]);
$fdisplay(file, "0x66A0,0x%h_0x%h", db_odd.mem_bank[821],db_even.mem_bank[821]);
$fdisplay(file, "0x66C0,0x%h_0x%h", db_odd.mem_bank[822],db_even.mem_bank[822]);
$fdisplay(file, "0x66E0,0x%h_0x%h", db_odd.mem_bank[823],db_even.mem_bank[823]);
$fdisplay(file, "0x6700,0x%h_0x%h", db_odd.mem_bank[824],db_even.mem_bank[824]);
$fdisplay(file, "0x6720,0x%h_0x%h", db_odd.mem_bank[825],db_even.mem_bank[825]);
$fdisplay(file, "0x6740,0x%h_0x%h", db_odd.mem_bank[826],db_even.mem_bank[826]);
$fdisplay(file, "0x6760,0x%h_0x%h", db_odd.mem_bank[827],db_even.mem_bank[827]);
$fdisplay(file, "0x6780,0x%h_0x%h", db_odd.mem_bank[828],db_even.mem_bank[828]);
$fdisplay(file, "0x67A0,0x%h_0x%h", db_odd.mem_bank[829],db_even.mem_bank[829]);
$fdisplay(file, "0x67C0,0x%h_0x%h", db_odd.mem_bank[830],db_even.mem_bank[830]);
$fdisplay(file, "0x67E0,0x%h_0x%h", db_odd.mem_bank[831],db_even.mem_bank[831]);
$fdisplay(file, "0x6800,0x%h_0x%h", db_odd.mem_bank[832],db_even.mem_bank[832]);
$fdisplay(file, "0x6820,0x%h_0x%h", db_odd.mem_bank[833],db_even.mem_bank[833]);
$fdisplay(file, "0x6840,0x%h_0x%h", db_odd.mem_bank[834],db_even.mem_bank[834]);
$fdisplay(file, "0x6860,0x%h_0x%h", db_odd.mem_bank[835],db_even.mem_bank[835]);
$fdisplay(file, "0x6880,0x%h_0x%h", db_odd.mem_bank[836],db_even.mem_bank[836]);
$fdisplay(file, "0x68A0,0x%h_0x%h", db_odd.mem_bank[837],db_even.mem_bank[837]);
$fdisplay(file, "0x68C0,0x%h_0x%h", db_odd.mem_bank[838],db_even.mem_bank[838]);
$fdisplay(file, "0x68E0,0x%h_0x%h", db_odd.mem_bank[839],db_even.mem_bank[839]);
$fdisplay(file, "0x6900,0x%h_0x%h", db_odd.mem_bank[840],db_even.mem_bank[840]);
$fdisplay(file, "0x6920,0x%h_0x%h", db_odd.mem_bank[841],db_even.mem_bank[841]);
$fdisplay(file, "0x6940,0x%h_0x%h", db_odd.mem_bank[842],db_even.mem_bank[842]);
$fdisplay(file, "0x6960,0x%h_0x%h", db_odd.mem_bank[843],db_even.mem_bank[843]);
$fdisplay(file, "0x6980,0x%h_0x%h", db_odd.mem_bank[844],db_even.mem_bank[844]);
$fdisplay(file, "0x69A0,0x%h_0x%h", db_odd.mem_bank[845],db_even.mem_bank[845]);
$fdisplay(file, "0x69C0,0x%h_0x%h", db_odd.mem_bank[846],db_even.mem_bank[846]);
$fdisplay(file, "0x69E0,0x%h_0x%h", db_odd.mem_bank[847],db_even.mem_bank[847]);
$fdisplay(file, "0x6A00,0x%h_0x%h", db_odd.mem_bank[848],db_even.mem_bank[848]);
$fdisplay(file, "0x6A20,0x%h_0x%h", db_odd.mem_bank[849],db_even.mem_bank[849]);
$fdisplay(file, "0x6A40,0x%h_0x%h", db_odd.mem_bank[850],db_even.mem_bank[850]);
$fdisplay(file, "0x6A60,0x%h_0x%h", db_odd.mem_bank[851],db_even.mem_bank[851]);
$fdisplay(file, "0x6A80,0x%h_0x%h", db_odd.mem_bank[852],db_even.mem_bank[852]);
$fdisplay(file, "0x6AA0,0x%h_0x%h", db_odd.mem_bank[853],db_even.mem_bank[853]);
$fdisplay(file, "0x6AC0,0x%h_0x%h", db_odd.mem_bank[854],db_even.mem_bank[854]);
$fdisplay(file, "0x6AE0,0x%h_0x%h", db_odd.mem_bank[855],db_even.mem_bank[855]);
$fdisplay(file, "0x6B00,0x%h_0x%h", db_odd.mem_bank[856],db_even.mem_bank[856]);
$fdisplay(file, "0x6B20,0x%h_0x%h", db_odd.mem_bank[857],db_even.mem_bank[857]);
$fdisplay(file, "0x6B40,0x%h_0x%h", db_odd.mem_bank[858],db_even.mem_bank[858]);
$fdisplay(file, "0x6B60,0x%h_0x%h", db_odd.mem_bank[859],db_even.mem_bank[859]);
$fdisplay(file, "0x6B80,0x%h_0x%h", db_odd.mem_bank[860],db_even.mem_bank[860]);
$fdisplay(file, "0x6BA0,0x%h_0x%h", db_odd.mem_bank[861],db_even.mem_bank[861]);
$fdisplay(file, "0x6BC0,0x%h_0x%h", db_odd.mem_bank[862],db_even.mem_bank[862]);
$fdisplay(file, "0x6BE0,0x%h_0x%h", db_odd.mem_bank[863],db_even.mem_bank[863]);
$fdisplay(file, "0x6C00,0x%h_0x%h", db_odd.mem_bank[864],db_even.mem_bank[864]);
$fdisplay(file, "0x6C20,0x%h_0x%h", db_odd.mem_bank[865],db_even.mem_bank[865]);
$fdisplay(file, "0x6C40,0x%h_0x%h", db_odd.mem_bank[866],db_even.mem_bank[866]);
$fdisplay(file, "0x6C60,0x%h_0x%h", db_odd.mem_bank[867],db_even.mem_bank[867]);
$fdisplay(file, "0x6C80,0x%h_0x%h", db_odd.mem_bank[868],db_even.mem_bank[868]);
$fdisplay(file, "0x6CA0,0x%h_0x%h", db_odd.mem_bank[869],db_even.mem_bank[869]);
$fdisplay(file, "0x6CC0,0x%h_0x%h", db_odd.mem_bank[870],db_even.mem_bank[870]);
$fdisplay(file, "0x6CE0,0x%h_0x%h", db_odd.mem_bank[871],db_even.mem_bank[871]);
$fdisplay(file, "0x6D00,0x%h_0x%h", db_odd.mem_bank[872],db_even.mem_bank[872]);
$fdisplay(file, "0x6D20,0x%h_0x%h", db_odd.mem_bank[873],db_even.mem_bank[873]);
$fdisplay(file, "0x6D40,0x%h_0x%h", db_odd.mem_bank[874],db_even.mem_bank[874]);
$fdisplay(file, "0x6D60,0x%h_0x%h", db_odd.mem_bank[875],db_even.mem_bank[875]);
$fdisplay(file, "0x6D80,0x%h_0x%h", db_odd.mem_bank[876],db_even.mem_bank[876]);
$fdisplay(file, "0x6DA0,0x%h_0x%h", db_odd.mem_bank[877],db_even.mem_bank[877]);
$fdisplay(file, "0x6DC0,0x%h_0x%h", db_odd.mem_bank[878],db_even.mem_bank[878]);
$fdisplay(file, "0x6DE0,0x%h_0x%h", db_odd.mem_bank[879],db_even.mem_bank[879]);
$fdisplay(file, "0x6E00,0x%h_0x%h", db_odd.mem_bank[880],db_even.mem_bank[880]);
$fdisplay(file, "0x6E20,0x%h_0x%h", db_odd.mem_bank[881],db_even.mem_bank[881]);
$fdisplay(file, "0x6E40,0x%h_0x%h", db_odd.mem_bank[882],db_even.mem_bank[882]);
$fdisplay(file, "0x6E60,0x%h_0x%h", db_odd.mem_bank[883],db_even.mem_bank[883]);
$fdisplay(file, "0x6E80,0x%h_0x%h", db_odd.mem_bank[884],db_even.mem_bank[884]);
$fdisplay(file, "0x6EA0,0x%h_0x%h", db_odd.mem_bank[885],db_even.mem_bank[885]);
$fdisplay(file, "0x6EC0,0x%h_0x%h", db_odd.mem_bank[886],db_even.mem_bank[886]);
$fdisplay(file, "0x6EE0,0x%h_0x%h", db_odd.mem_bank[887],db_even.mem_bank[887]);
$fdisplay(file, "0x6F00,0x%h_0x%h", db_odd.mem_bank[888],db_even.mem_bank[888]);
$fdisplay(file, "0x6F20,0x%h_0x%h", db_odd.mem_bank[889],db_even.mem_bank[889]);
$fdisplay(file, "0x6F40,0x%h_0x%h", db_odd.mem_bank[890],db_even.mem_bank[890]);
$fdisplay(file, "0x6F60,0x%h_0x%h", db_odd.mem_bank[891],db_even.mem_bank[891]);
$fdisplay(file, "0x6F80,0x%h_0x%h", db_odd.mem_bank[892],db_even.mem_bank[892]);
$fdisplay(file, "0x6FA0,0x%h_0x%h", db_odd.mem_bank[893],db_even.mem_bank[893]);
$fdisplay(file, "0x6FC0,0x%h_0x%h", db_odd.mem_bank[894],db_even.mem_bank[894]);
$fdisplay(file, "0x6FE0,0x%h_0x%h", db_odd.mem_bank[895],db_even.mem_bank[895]);
$fdisplay(file, "0x7000,0x%h_0x%h", db_odd.mem_bank[896],db_even.mem_bank[896]);
$fdisplay(file, "0x7020,0x%h_0x%h", db_odd.mem_bank[897],db_even.mem_bank[897]);
$fdisplay(file, "0x7040,0x%h_0x%h", db_odd.mem_bank[898],db_even.mem_bank[898]);
$fdisplay(file, "0x7060,0x%h_0x%h", db_odd.mem_bank[899],db_even.mem_bank[899]);
$fdisplay(file, "0x7080,0x%h_0x%h", db_odd.mem_bank[900],db_even.mem_bank[900]);
$fdisplay(file, "0x70A0,0x%h_0x%h", db_odd.mem_bank[901],db_even.mem_bank[901]);
$fdisplay(file, "0x70C0,0x%h_0x%h", db_odd.mem_bank[902],db_even.mem_bank[902]);
$fdisplay(file, "0x70E0,0x%h_0x%h", db_odd.mem_bank[903],db_even.mem_bank[903]);
$fdisplay(file, "0x7100,0x%h_0x%h", db_odd.mem_bank[904],db_even.mem_bank[904]);
$fdisplay(file, "0x7120,0x%h_0x%h", db_odd.mem_bank[905],db_even.mem_bank[905]);
$fdisplay(file, "0x7140,0x%h_0x%h", db_odd.mem_bank[906],db_even.mem_bank[906]);
$fdisplay(file, "0x7160,0x%h_0x%h", db_odd.mem_bank[907],db_even.mem_bank[907]);
$fdisplay(file, "0x7180,0x%h_0x%h", db_odd.mem_bank[908],db_even.mem_bank[908]);
$fdisplay(file, "0x71A0,0x%h_0x%h", db_odd.mem_bank[909],db_even.mem_bank[909]);
$fdisplay(file, "0x71C0,0x%h_0x%h", db_odd.mem_bank[910],db_even.mem_bank[910]);
$fdisplay(file, "0x71E0,0x%h_0x%h", db_odd.mem_bank[911],db_even.mem_bank[911]);
$fdisplay(file, "0x7200,0x%h_0x%h", db_odd.mem_bank[912],db_even.mem_bank[912]);
$fdisplay(file, "0x7220,0x%h_0x%h", db_odd.mem_bank[913],db_even.mem_bank[913]);
$fdisplay(file, "0x7240,0x%h_0x%h", db_odd.mem_bank[914],db_even.mem_bank[914]);
$fdisplay(file, "0x7260,0x%h_0x%h", db_odd.mem_bank[915],db_even.mem_bank[915]);
$fdisplay(file, "0x7280,0x%h_0x%h", db_odd.mem_bank[916],db_even.mem_bank[916]);
$fdisplay(file, "0x72A0,0x%h_0x%h", db_odd.mem_bank[917],db_even.mem_bank[917]);
$fdisplay(file, "0x72C0,0x%h_0x%h", db_odd.mem_bank[918],db_even.mem_bank[918]);
$fdisplay(file, "0x72E0,0x%h_0x%h", db_odd.mem_bank[919],db_even.mem_bank[919]);
$fdisplay(file, "0x7300,0x%h_0x%h", db_odd.mem_bank[920],db_even.mem_bank[920]);
$fdisplay(file, "0x7320,0x%h_0x%h", db_odd.mem_bank[921],db_even.mem_bank[921]);
$fdisplay(file, "0x7340,0x%h_0x%h", db_odd.mem_bank[922],db_even.mem_bank[922]);
$fdisplay(file, "0x7360,0x%h_0x%h", db_odd.mem_bank[923],db_even.mem_bank[923]);
$fdisplay(file, "0x7380,0x%h_0x%h", db_odd.mem_bank[924],db_even.mem_bank[924]);
$fdisplay(file, "0x73A0,0x%h_0x%h", db_odd.mem_bank[925],db_even.mem_bank[925]);
$fdisplay(file, "0x73C0,0x%h_0x%h", db_odd.mem_bank[926],db_even.mem_bank[926]);
$fdisplay(file, "0x73E0,0x%h_0x%h", db_odd.mem_bank[927],db_even.mem_bank[927]);
$fdisplay(file, "0x7400,0x%h_0x%h", db_odd.mem_bank[928],db_even.mem_bank[928]);
$fdisplay(file, "0x7420,0x%h_0x%h", db_odd.mem_bank[929],db_even.mem_bank[929]);
$fdisplay(file, "0x7440,0x%h_0x%h", db_odd.mem_bank[930],db_even.mem_bank[930]);
$fdisplay(file, "0x7460,0x%h_0x%h", db_odd.mem_bank[931],db_even.mem_bank[931]);
$fdisplay(file, "0x7480,0x%h_0x%h", db_odd.mem_bank[932],db_even.mem_bank[932]);
$fdisplay(file, "0x74A0,0x%h_0x%h", db_odd.mem_bank[933],db_even.mem_bank[933]);
$fdisplay(file, "0x74C0,0x%h_0x%h", db_odd.mem_bank[934],db_even.mem_bank[934]);
$fdisplay(file, "0x74E0,0x%h_0x%h", db_odd.mem_bank[935],db_even.mem_bank[935]);
$fdisplay(file, "0x7500,0x%h_0x%h", db_odd.mem_bank[936],db_even.mem_bank[936]);
$fdisplay(file, "0x7520,0x%h_0x%h", db_odd.mem_bank[937],db_even.mem_bank[937]);
$fdisplay(file, "0x7540,0x%h_0x%h", db_odd.mem_bank[938],db_even.mem_bank[938]);
$fdisplay(file, "0x7560,0x%h_0x%h", db_odd.mem_bank[939],db_even.mem_bank[939]);
$fdisplay(file, "0x7580,0x%h_0x%h", db_odd.mem_bank[940],db_even.mem_bank[940]);
$fdisplay(file, "0x75A0,0x%h_0x%h", db_odd.mem_bank[941],db_even.mem_bank[941]);
$fdisplay(file, "0x75C0,0x%h_0x%h", db_odd.mem_bank[942],db_even.mem_bank[942]);
$fdisplay(file, "0x75E0,0x%h_0x%h", db_odd.mem_bank[943],db_even.mem_bank[943]);
$fdisplay(file, "0x7600,0x%h_0x%h", db_odd.mem_bank[944],db_even.mem_bank[944]);
$fdisplay(file, "0x7620,0x%h_0x%h", db_odd.mem_bank[945],db_even.mem_bank[945]);
$fdisplay(file, "0x7640,0x%h_0x%h", db_odd.mem_bank[946],db_even.mem_bank[946]);
$fdisplay(file, "0x7660,0x%h_0x%h", db_odd.mem_bank[947],db_even.mem_bank[947]);
$fdisplay(file, "0x7680,0x%h_0x%h", db_odd.mem_bank[948],db_even.mem_bank[948]);
$fdisplay(file, "0x76A0,0x%h_0x%h", db_odd.mem_bank[949],db_even.mem_bank[949]);
$fdisplay(file, "0x76C0,0x%h_0x%h", db_odd.mem_bank[950],db_even.mem_bank[950]);
$fdisplay(file, "0x76E0,0x%h_0x%h", db_odd.mem_bank[951],db_even.mem_bank[951]);
$fdisplay(file, "0x7700,0x%h_0x%h", db_odd.mem_bank[952],db_even.mem_bank[952]);
$fdisplay(file, "0x7720,0x%h_0x%h", db_odd.mem_bank[953],db_even.mem_bank[953]);
$fdisplay(file, "0x7740,0x%h_0x%h", db_odd.mem_bank[954],db_even.mem_bank[954]);
$fdisplay(file, "0x7760,0x%h_0x%h", db_odd.mem_bank[955],db_even.mem_bank[955]);
$fdisplay(file, "0x7780,0x%h_0x%h", db_odd.mem_bank[956],db_even.mem_bank[956]);
$fdisplay(file, "0x77A0,0x%h_0x%h", db_odd.mem_bank[957],db_even.mem_bank[957]);
$fdisplay(file, "0x77C0,0x%h_0x%h", db_odd.mem_bank[958],db_even.mem_bank[958]);
$fdisplay(file, "0x77E0,0x%h_0x%h", db_odd.mem_bank[959],db_even.mem_bank[959]);
$fdisplay(file, "0x7800,0x%h_0x%h", db_odd.mem_bank[960],db_even.mem_bank[960]);
$fdisplay(file, "0x7820,0x%h_0x%h", db_odd.mem_bank[961],db_even.mem_bank[961]);
$fdisplay(file, "0x7840,0x%h_0x%h", db_odd.mem_bank[962],db_even.mem_bank[962]);
$fdisplay(file, "0x7860,0x%h_0x%h", db_odd.mem_bank[963],db_even.mem_bank[963]);
$fdisplay(file, "0x7880,0x%h_0x%h", db_odd.mem_bank[964],db_even.mem_bank[964]);
$fdisplay(file, "0x78A0,0x%h_0x%h", db_odd.mem_bank[965],db_even.mem_bank[965]);
$fdisplay(file, "0x78C0,0x%h_0x%h", db_odd.mem_bank[966],db_even.mem_bank[966]);
$fdisplay(file, "0x78E0,0x%h_0x%h", db_odd.mem_bank[967],db_even.mem_bank[967]);
$fdisplay(file, "0x7900,0x%h_0x%h", db_odd.mem_bank[968],db_even.mem_bank[968]);
$fdisplay(file, "0x7920,0x%h_0x%h", db_odd.mem_bank[969],db_even.mem_bank[969]);
$fdisplay(file, "0x7940,0x%h_0x%h", db_odd.mem_bank[970],db_even.mem_bank[970]);
$fdisplay(file, "0x7960,0x%h_0x%h", db_odd.mem_bank[971],db_even.mem_bank[971]);
$fdisplay(file, "0x7980,0x%h_0x%h", db_odd.mem_bank[972],db_even.mem_bank[972]);
$fdisplay(file, "0x79A0,0x%h_0x%h", db_odd.mem_bank[973],db_even.mem_bank[973]);
$fdisplay(file, "0x79C0,0x%h_0x%h", db_odd.mem_bank[974],db_even.mem_bank[974]);
$fdisplay(file, "0x79E0,0x%h_0x%h", db_odd.mem_bank[975],db_even.mem_bank[975]);
$fdisplay(file, "0x7A00,0x%h_0x%h", db_odd.mem_bank[976],db_even.mem_bank[976]);
$fdisplay(file, "0x7A20,0x%h_0x%h", db_odd.mem_bank[977],db_even.mem_bank[977]);
$fdisplay(file, "0x7A40,0x%h_0x%h", db_odd.mem_bank[978],db_even.mem_bank[978]);
$fdisplay(file, "0x7A60,0x%h_0x%h", db_odd.mem_bank[979],db_even.mem_bank[979]);
$fdisplay(file, "0x7A80,0x%h_0x%h", db_odd.mem_bank[980],db_even.mem_bank[980]);
$fdisplay(file, "0x7AA0,0x%h_0x%h", db_odd.mem_bank[981],db_even.mem_bank[981]);
$fdisplay(file, "0x7AC0,0x%h_0x%h", db_odd.mem_bank[982],db_even.mem_bank[982]);
$fdisplay(file, "0x7AE0,0x%h_0x%h", db_odd.mem_bank[983],db_even.mem_bank[983]);
$fdisplay(file, "0x7B00,0x%h_0x%h", db_odd.mem_bank[984],db_even.mem_bank[984]);
$fdisplay(file, "0x7B20,0x%h_0x%h", db_odd.mem_bank[985],db_even.mem_bank[985]);
$fdisplay(file, "0x7B40,0x%h_0x%h", db_odd.mem_bank[986],db_even.mem_bank[986]);
$fdisplay(file, "0x7B60,0x%h_0x%h", db_odd.mem_bank[987],db_even.mem_bank[987]);
$fdisplay(file, "0x7B80,0x%h_0x%h", db_odd.mem_bank[988],db_even.mem_bank[988]);
$fdisplay(file, "0x7BA0,0x%h_0x%h", db_odd.mem_bank[989],db_even.mem_bank[989]);
$fdisplay(file, "0x7BC0,0x%h_0x%h", db_odd.mem_bank[990],db_even.mem_bank[990]);
$fdisplay(file, "0x7BE0,0x%h_0x%h", db_odd.mem_bank[991],db_even.mem_bank[991]);
$fdisplay(file, "0x7C00,0x%h_0x%h", db_odd.mem_bank[992],db_even.mem_bank[992]);
$fdisplay(file, "0x7C20,0x%h_0x%h", db_odd.mem_bank[993],db_even.mem_bank[993]);
$fdisplay(file, "0x7C40,0x%h_0x%h", db_odd.mem_bank[994],db_even.mem_bank[994]);
$fdisplay(file, "0x7C60,0x%h_0x%h", db_odd.mem_bank[995],db_even.mem_bank[995]);
$fdisplay(file, "0x7C80,0x%h_0x%h", db_odd.mem_bank[996],db_even.mem_bank[996]);
$fdisplay(file, "0x7CA0,0x%h_0x%h", db_odd.mem_bank[997],db_even.mem_bank[997]);
$fdisplay(file, "0x7CC0,0x%h_0x%h", db_odd.mem_bank[998],db_even.mem_bank[998]);
$fdisplay(file, "0x7CE0,0x%h_0x%h", db_odd.mem_bank[999],db_even.mem_bank[999]);
$fdisplay(file, "0x7D00,0x%h_0x%h", db_odd.mem_bank[1000],db_even.mem_bank[1000]);
$fdisplay(file, "0x7D20,0x%h_0x%h", db_odd.mem_bank[1001],db_even.mem_bank[1001]);
$fdisplay(file, "0x7D40,0x%h_0x%h", db_odd.mem_bank[1002],db_even.mem_bank[1002]);
$fdisplay(file, "0x7D60,0x%h_0x%h", db_odd.mem_bank[1003],db_even.mem_bank[1003]);
$fdisplay(file, "0x7D80,0x%h_0x%h", db_odd.mem_bank[1004],db_even.mem_bank[1004]);
$fdisplay(file, "0x7DA0,0x%h_0x%h", db_odd.mem_bank[1005],db_even.mem_bank[1005]);
$fdisplay(file, "0x7DC0,0x%h_0x%h", db_odd.mem_bank[1006],db_even.mem_bank[1006]);
$fdisplay(file, "0x7DE0,0x%h_0x%h", db_odd.mem_bank[1007],db_even.mem_bank[1007]);
$fdisplay(file, "0x7E00,0x%h_0x%h", db_odd.mem_bank[1008],db_even.mem_bank[1008]);
$fdisplay(file, "0x7E20,0x%h_0x%h", db_odd.mem_bank[1009],db_even.mem_bank[1009]);
$fdisplay(file, "0x7E40,0x%h_0x%h", db_odd.mem_bank[1010],db_even.mem_bank[1010]);
$fdisplay(file, "0x7E60,0x%h_0x%h", db_odd.mem_bank[1011],db_even.mem_bank[1011]);
$fdisplay(file, "0x7E80,0x%h_0x%h", db_odd.mem_bank[1012],db_even.mem_bank[1012]);
$fdisplay(file, "0x7EA0,0x%h_0x%h", db_odd.mem_bank[1013],db_even.mem_bank[1013]);
$fdisplay(file, "0x7EC0,0x%h_0x%h", db_odd.mem_bank[1014],db_even.mem_bank[1014]);
$fdisplay(file, "0x7EE0,0x%h_0x%h", db_odd.mem_bank[1015],db_even.mem_bank[1015]);
$fdisplay(file, "0x7F00,0x%h_0x%h", db_odd.mem_bank[1016],db_even.mem_bank[1016]);
$fdisplay(file, "0x7F20,0x%h_0x%h", db_odd.mem_bank[1017],db_even.mem_bank[1017]);
$fdisplay(file, "0x7F40,0x%h_0x%h", db_odd.mem_bank[1018],db_even.mem_bank[1018]);
$fdisplay(file, "0x7F60,0x%h_0x%h", db_odd.mem_bank[1019],db_even.mem_bank[1019]);
$fdisplay(file, "0x7F80,0x%h_0x%h", db_odd.mem_bank[1020],db_even.mem_bank[1020]);
$fdisplay(file, "0x7FA0,0x%h_0x%h", db_odd.mem_bank[1021],db_even.mem_bank[1021]);
$fdisplay(file, "0x7FC0,0x%h_0x%h", db_odd.mem_bank[1022],db_even.mem_bank[1022]);
$fdisplay(file, "0x7FE0,0x%h_0x%h", db_odd.mem_bank[1023],db_even.mem_bank[1023]);
$fdisplay(file, "0x8000,0x%h_0x%h", db_odd.mem_bank[1024],db_even.mem_bank[1024]);
$fdisplay(file, "0x8020,0x%h_0x%h", db_odd.mem_bank[1025],db_even.mem_bank[1025]);
$fdisplay(file, "0x8040,0x%h_0x%h", db_odd.mem_bank[1026],db_even.mem_bank[1026]);
$fdisplay(file, "0x8060,0x%h_0x%h", db_odd.mem_bank[1027],db_even.mem_bank[1027]);
$fdisplay(file, "0x8080,0x%h_0x%h", db_odd.mem_bank[1028],db_even.mem_bank[1028]);
$fdisplay(file, "0x80A0,0x%h_0x%h", db_odd.mem_bank[1029],db_even.mem_bank[1029]);
$fdisplay(file, "0x80C0,0x%h_0x%h", db_odd.mem_bank[1030],db_even.mem_bank[1030]);
$fdisplay(file, "0x80E0,0x%h_0x%h", db_odd.mem_bank[1031],db_even.mem_bank[1031]);
$fdisplay(file, "0x8100,0x%h_0x%h", db_odd.mem_bank[1032],db_even.mem_bank[1032]);
$fdisplay(file, "0x8120,0x%h_0x%h", db_odd.mem_bank[1033],db_even.mem_bank[1033]);
$fdisplay(file, "0x8140,0x%h_0x%h", db_odd.mem_bank[1034],db_even.mem_bank[1034]);
$fdisplay(file, "0x8160,0x%h_0x%h", db_odd.mem_bank[1035],db_even.mem_bank[1035]);
$fdisplay(file, "0x8180,0x%h_0x%h", db_odd.mem_bank[1036],db_even.mem_bank[1036]);
$fdisplay(file, "0x81A0,0x%h_0x%h", db_odd.mem_bank[1037],db_even.mem_bank[1037]);
$fdisplay(file, "0x81C0,0x%h_0x%h", db_odd.mem_bank[1038],db_even.mem_bank[1038]);
$fdisplay(file, "0x81E0,0x%h_0x%h", db_odd.mem_bank[1039],db_even.mem_bank[1039]);
$fdisplay(file, "0x8200,0x%h_0x%h", db_odd.mem_bank[1040],db_even.mem_bank[1040]);
$fdisplay(file, "0x8220,0x%h_0x%h", db_odd.mem_bank[1041],db_even.mem_bank[1041]);
$fdisplay(file, "0x8240,0x%h_0x%h", db_odd.mem_bank[1042],db_even.mem_bank[1042]);
$fdisplay(file, "0x8260,0x%h_0x%h", db_odd.mem_bank[1043],db_even.mem_bank[1043]);
$fdisplay(file, "0x8280,0x%h_0x%h", db_odd.mem_bank[1044],db_even.mem_bank[1044]);
$fdisplay(file, "0x82A0,0x%h_0x%h", db_odd.mem_bank[1045],db_even.mem_bank[1045]);
$fdisplay(file, "0x82C0,0x%h_0x%h", db_odd.mem_bank[1046],db_even.mem_bank[1046]);
$fdisplay(file, "0x82E0,0x%h_0x%h", db_odd.mem_bank[1047],db_even.mem_bank[1047]);
$fdisplay(file, "0x8300,0x%h_0x%h", db_odd.mem_bank[1048],db_even.mem_bank[1048]);
$fdisplay(file, "0x8320,0x%h_0x%h", db_odd.mem_bank[1049],db_even.mem_bank[1049]);
$fdisplay(file, "0x8340,0x%h_0x%h", db_odd.mem_bank[1050],db_even.mem_bank[1050]);
$fdisplay(file, "0x8360,0x%h_0x%h", db_odd.mem_bank[1051],db_even.mem_bank[1051]);
$fdisplay(file, "0x8380,0x%h_0x%h", db_odd.mem_bank[1052],db_even.mem_bank[1052]);
$fdisplay(file, "0x83A0,0x%h_0x%h", db_odd.mem_bank[1053],db_even.mem_bank[1053]);
$fdisplay(file, "0x83C0,0x%h_0x%h", db_odd.mem_bank[1054],db_even.mem_bank[1054]);
$fdisplay(file, "0x83E0,0x%h_0x%h", db_odd.mem_bank[1055],db_even.mem_bank[1055]);
$fdisplay(file, "0x8400,0x%h_0x%h", db_odd.mem_bank[1056],db_even.mem_bank[1056]);
$fdisplay(file, "0x8420,0x%h_0x%h", db_odd.mem_bank[1057],db_even.mem_bank[1057]);
$fdisplay(file, "0x8440,0x%h_0x%h", db_odd.mem_bank[1058],db_even.mem_bank[1058]);
$fdisplay(file, "0x8460,0x%h_0x%h", db_odd.mem_bank[1059],db_even.mem_bank[1059]);
$fdisplay(file, "0x8480,0x%h_0x%h", db_odd.mem_bank[1060],db_even.mem_bank[1060]);
$fdisplay(file, "0x84A0,0x%h_0x%h", db_odd.mem_bank[1061],db_even.mem_bank[1061]);
$fdisplay(file, "0x84C0,0x%h_0x%h", db_odd.mem_bank[1062],db_even.mem_bank[1062]);
$fdisplay(file, "0x84E0,0x%h_0x%h", db_odd.mem_bank[1063],db_even.mem_bank[1063]);
$fdisplay(file, "0x8500,0x%h_0x%h", db_odd.mem_bank[1064],db_even.mem_bank[1064]);
$fdisplay(file, "0x8520,0x%h_0x%h", db_odd.mem_bank[1065],db_even.mem_bank[1065]);
$fdisplay(file, "0x8540,0x%h_0x%h", db_odd.mem_bank[1066],db_even.mem_bank[1066]);
$fdisplay(file, "0x8560,0x%h_0x%h", db_odd.mem_bank[1067],db_even.mem_bank[1067]);
$fdisplay(file, "0x8580,0x%h_0x%h", db_odd.mem_bank[1068],db_even.mem_bank[1068]);
$fdisplay(file, "0x85A0,0x%h_0x%h", db_odd.mem_bank[1069],db_even.mem_bank[1069]);
$fdisplay(file, "0x85C0,0x%h_0x%h", db_odd.mem_bank[1070],db_even.mem_bank[1070]);
$fdisplay(file, "0x85E0,0x%h_0x%h", db_odd.mem_bank[1071],db_even.mem_bank[1071]);
$fdisplay(file, "0x8600,0x%h_0x%h", db_odd.mem_bank[1072],db_even.mem_bank[1072]);
$fdisplay(file, "0x8620,0x%h_0x%h", db_odd.mem_bank[1073],db_even.mem_bank[1073]);
$fdisplay(file, "0x8640,0x%h_0x%h", db_odd.mem_bank[1074],db_even.mem_bank[1074]);
$fdisplay(file, "0x8660,0x%h_0x%h", db_odd.mem_bank[1075],db_even.mem_bank[1075]);
$fdisplay(file, "0x8680,0x%h_0x%h", db_odd.mem_bank[1076],db_even.mem_bank[1076]);
$fdisplay(file, "0x86A0,0x%h_0x%h", db_odd.mem_bank[1077],db_even.mem_bank[1077]);
$fdisplay(file, "0x86C0,0x%h_0x%h", db_odd.mem_bank[1078],db_even.mem_bank[1078]);
$fdisplay(file, "0x86E0,0x%h_0x%h", db_odd.mem_bank[1079],db_even.mem_bank[1079]);
$fdisplay(file, "0x8700,0x%h_0x%h", db_odd.mem_bank[1080],db_even.mem_bank[1080]);
$fdisplay(file, "0x8720,0x%h_0x%h", db_odd.mem_bank[1081],db_even.mem_bank[1081]);
$fdisplay(file, "0x8740,0x%h_0x%h", db_odd.mem_bank[1082],db_even.mem_bank[1082]);
$fdisplay(file, "0x8760,0x%h_0x%h", db_odd.mem_bank[1083],db_even.mem_bank[1083]);
$fdisplay(file, "0x8780,0x%h_0x%h", db_odd.mem_bank[1084],db_even.mem_bank[1084]);
$fdisplay(file, "0x87A0,0x%h_0x%h", db_odd.mem_bank[1085],db_even.mem_bank[1085]);
$fdisplay(file, "0x87C0,0x%h_0x%h", db_odd.mem_bank[1086],db_even.mem_bank[1086]);
$fdisplay(file, "0x87E0,0x%h_0x%h", db_odd.mem_bank[1087],db_even.mem_bank[1087]);
$fdisplay(file, "0x8800,0x%h_0x%h", db_odd.mem_bank[1088],db_even.mem_bank[1088]);
$fdisplay(file, "0x8820,0x%h_0x%h", db_odd.mem_bank[1089],db_even.mem_bank[1089]);
$fdisplay(file, "0x8840,0x%h_0x%h", db_odd.mem_bank[1090],db_even.mem_bank[1090]);
$fdisplay(file, "0x8860,0x%h_0x%h", db_odd.mem_bank[1091],db_even.mem_bank[1091]);
$fdisplay(file, "0x8880,0x%h_0x%h", db_odd.mem_bank[1092],db_even.mem_bank[1092]);
$fdisplay(file, "0x88A0,0x%h_0x%h", db_odd.mem_bank[1093],db_even.mem_bank[1093]);
$fdisplay(file, "0x88C0,0x%h_0x%h", db_odd.mem_bank[1094],db_even.mem_bank[1094]);
$fdisplay(file, "0x88E0,0x%h_0x%h", db_odd.mem_bank[1095],db_even.mem_bank[1095]);
$fdisplay(file, "0x8900,0x%h_0x%h", db_odd.mem_bank[1096],db_even.mem_bank[1096]);
$fdisplay(file, "0x8920,0x%h_0x%h", db_odd.mem_bank[1097],db_even.mem_bank[1097]);
$fdisplay(file, "0x8940,0x%h_0x%h", db_odd.mem_bank[1098],db_even.mem_bank[1098]);
$fdisplay(file, "0x8960,0x%h_0x%h", db_odd.mem_bank[1099],db_even.mem_bank[1099]);
$fdisplay(file, "0x8980,0x%h_0x%h", db_odd.mem_bank[1100],db_even.mem_bank[1100]);
$fdisplay(file, "0x89A0,0x%h_0x%h", db_odd.mem_bank[1101],db_even.mem_bank[1101]);
$fdisplay(file, "0x89C0,0x%h_0x%h", db_odd.mem_bank[1102],db_even.mem_bank[1102]);
$fdisplay(file, "0x89E0,0x%h_0x%h", db_odd.mem_bank[1103],db_even.mem_bank[1103]);
$fdisplay(file, "0x8A00,0x%h_0x%h", db_odd.mem_bank[1104],db_even.mem_bank[1104]);
$fdisplay(file, "0x8A20,0x%h_0x%h", db_odd.mem_bank[1105],db_even.mem_bank[1105]);
$fdisplay(file, "0x8A40,0x%h_0x%h", db_odd.mem_bank[1106],db_even.mem_bank[1106]);
$fdisplay(file, "0x8A60,0x%h_0x%h", db_odd.mem_bank[1107],db_even.mem_bank[1107]);
$fdisplay(file, "0x8A80,0x%h_0x%h", db_odd.mem_bank[1108],db_even.mem_bank[1108]);
$fdisplay(file, "0x8AA0,0x%h_0x%h", db_odd.mem_bank[1109],db_even.mem_bank[1109]);
$fdisplay(file, "0x8AC0,0x%h_0x%h", db_odd.mem_bank[1110],db_even.mem_bank[1110]);
$fdisplay(file, "0x8AE0,0x%h_0x%h", db_odd.mem_bank[1111],db_even.mem_bank[1111]);
$fdisplay(file, "0x8B00,0x%h_0x%h", db_odd.mem_bank[1112],db_even.mem_bank[1112]);
$fdisplay(file, "0x8B20,0x%h_0x%h", db_odd.mem_bank[1113],db_even.mem_bank[1113]);
$fdisplay(file, "0x8B40,0x%h_0x%h", db_odd.mem_bank[1114],db_even.mem_bank[1114]);
$fdisplay(file, "0x8B60,0x%h_0x%h", db_odd.mem_bank[1115],db_even.mem_bank[1115]);
$fdisplay(file, "0x8B80,0x%h_0x%h", db_odd.mem_bank[1116],db_even.mem_bank[1116]);
$fdisplay(file, "0x8BA0,0x%h_0x%h", db_odd.mem_bank[1117],db_even.mem_bank[1117]);
$fdisplay(file, "0x8BC0,0x%h_0x%h", db_odd.mem_bank[1118],db_even.mem_bank[1118]);
$fdisplay(file, "0x8BE0,0x%h_0x%h", db_odd.mem_bank[1119],db_even.mem_bank[1119]);
$fdisplay(file, "0x8C00,0x%h_0x%h", db_odd.mem_bank[1120],db_even.mem_bank[1120]);
$fdisplay(file, "0x8C20,0x%h_0x%h", db_odd.mem_bank[1121],db_even.mem_bank[1121]);
$fdisplay(file, "0x8C40,0x%h_0x%h", db_odd.mem_bank[1122],db_even.mem_bank[1122]);
$fdisplay(file, "0x8C60,0x%h_0x%h", db_odd.mem_bank[1123],db_even.mem_bank[1123]);
$fdisplay(file, "0x8C80,0x%h_0x%h", db_odd.mem_bank[1124],db_even.mem_bank[1124]);
$fdisplay(file, "0x8CA0,0x%h_0x%h", db_odd.mem_bank[1125],db_even.mem_bank[1125]);
$fdisplay(file, "0x8CC0,0x%h_0x%h", db_odd.mem_bank[1126],db_even.mem_bank[1126]);
$fdisplay(file, "0x8CE0,0x%h_0x%h", db_odd.mem_bank[1127],db_even.mem_bank[1127]);
$fdisplay(file, "0x8D00,0x%h_0x%h", db_odd.mem_bank[1128],db_even.mem_bank[1128]);
$fdisplay(file, "0x8D20,0x%h_0x%h", db_odd.mem_bank[1129],db_even.mem_bank[1129]);
$fdisplay(file, "0x8D40,0x%h_0x%h", db_odd.mem_bank[1130],db_even.mem_bank[1130]);
$fdisplay(file, "0x8D60,0x%h_0x%h", db_odd.mem_bank[1131],db_even.mem_bank[1131]);
$fdisplay(file, "0x8D80,0x%h_0x%h", db_odd.mem_bank[1132],db_even.mem_bank[1132]);
$fdisplay(file, "0x8DA0,0x%h_0x%h", db_odd.mem_bank[1133],db_even.mem_bank[1133]);
$fdisplay(file, "0x8DC0,0x%h_0x%h", db_odd.mem_bank[1134],db_even.mem_bank[1134]);
$fdisplay(file, "0x8DE0,0x%h_0x%h", db_odd.mem_bank[1135],db_even.mem_bank[1135]);
$fdisplay(file, "0x8E00,0x%h_0x%h", db_odd.mem_bank[1136],db_even.mem_bank[1136]);
$fdisplay(file, "0x8E20,0x%h_0x%h", db_odd.mem_bank[1137],db_even.mem_bank[1137]);
$fdisplay(file, "0x8E40,0x%h_0x%h", db_odd.mem_bank[1138],db_even.mem_bank[1138]);
$fdisplay(file, "0x8E60,0x%h_0x%h", db_odd.mem_bank[1139],db_even.mem_bank[1139]);
$fdisplay(file, "0x8E80,0x%h_0x%h", db_odd.mem_bank[1140],db_even.mem_bank[1140]);
$fdisplay(file, "0x8EA0,0x%h_0x%h", db_odd.mem_bank[1141],db_even.mem_bank[1141]);
$fdisplay(file, "0x8EC0,0x%h_0x%h", db_odd.mem_bank[1142],db_even.mem_bank[1142]);
$fdisplay(file, "0x8EE0,0x%h_0x%h", db_odd.mem_bank[1143],db_even.mem_bank[1143]);
$fdisplay(file, "0x8F00,0x%h_0x%h", db_odd.mem_bank[1144],db_even.mem_bank[1144]);
$fdisplay(file, "0x8F20,0x%h_0x%h", db_odd.mem_bank[1145],db_even.mem_bank[1145]);
$fdisplay(file, "0x8F40,0x%h_0x%h", db_odd.mem_bank[1146],db_even.mem_bank[1146]);
$fdisplay(file, "0x8F60,0x%h_0x%h", db_odd.mem_bank[1147],db_even.mem_bank[1147]);
$fdisplay(file, "0x8F80,0x%h_0x%h", db_odd.mem_bank[1148],db_even.mem_bank[1148]);
$fdisplay(file, "0x8FA0,0x%h_0x%h", db_odd.mem_bank[1149],db_even.mem_bank[1149]);
$fdisplay(file, "0x8FC0,0x%h_0x%h", db_odd.mem_bank[1150],db_even.mem_bank[1150]);
$fdisplay(file, "0x8FE0,0x%h_0x%h", db_odd.mem_bank[1151],db_even.mem_bank[1151]);
$fdisplay(file, "0x9000,0x%h_0x%h", db_odd.mem_bank[1152],db_even.mem_bank[1152]);
$fdisplay(file, "0x9020,0x%h_0x%h", db_odd.mem_bank[1153],db_even.mem_bank[1153]);
$fdisplay(file, "0x9040,0x%h_0x%h", db_odd.mem_bank[1154],db_even.mem_bank[1154]);
$fdisplay(file, "0x9060,0x%h_0x%h", db_odd.mem_bank[1155],db_even.mem_bank[1155]);
$fdisplay(file, "0x9080,0x%h_0x%h", db_odd.mem_bank[1156],db_even.mem_bank[1156]);
$fdisplay(file, "0x90A0,0x%h_0x%h", db_odd.mem_bank[1157],db_even.mem_bank[1157]);
$fdisplay(file, "0x90C0,0x%h_0x%h", db_odd.mem_bank[1158],db_even.mem_bank[1158]);
$fdisplay(file, "0x90E0,0x%h_0x%h", db_odd.mem_bank[1159],db_even.mem_bank[1159]);
$fdisplay(file, "0x9100,0x%h_0x%h", db_odd.mem_bank[1160],db_even.mem_bank[1160]);
$fdisplay(file, "0x9120,0x%h_0x%h", db_odd.mem_bank[1161],db_even.mem_bank[1161]);
$fdisplay(file, "0x9140,0x%h_0x%h", db_odd.mem_bank[1162],db_even.mem_bank[1162]);
$fdisplay(file, "0x9160,0x%h_0x%h", db_odd.mem_bank[1163],db_even.mem_bank[1163]);
$fdisplay(file, "0x9180,0x%h_0x%h", db_odd.mem_bank[1164],db_even.mem_bank[1164]);
$fdisplay(file, "0x91A0,0x%h_0x%h", db_odd.mem_bank[1165],db_even.mem_bank[1165]);
$fdisplay(file, "0x91C0,0x%h_0x%h", db_odd.mem_bank[1166],db_even.mem_bank[1166]);
$fdisplay(file, "0x91E0,0x%h_0x%h", db_odd.mem_bank[1167],db_even.mem_bank[1167]);
$fdisplay(file, "0x9200,0x%h_0x%h", db_odd.mem_bank[1168],db_even.mem_bank[1168]);
$fdisplay(file, "0x9220,0x%h_0x%h", db_odd.mem_bank[1169],db_even.mem_bank[1169]);
$fdisplay(file, "0x9240,0x%h_0x%h", db_odd.mem_bank[1170],db_even.mem_bank[1170]);
$fdisplay(file, "0x9260,0x%h_0x%h", db_odd.mem_bank[1171],db_even.mem_bank[1171]);
$fdisplay(file, "0x9280,0x%h_0x%h", db_odd.mem_bank[1172],db_even.mem_bank[1172]);
$fdisplay(file, "0x92A0,0x%h_0x%h", db_odd.mem_bank[1173],db_even.mem_bank[1173]);
$fdisplay(file, "0x92C0,0x%h_0x%h", db_odd.mem_bank[1174],db_even.mem_bank[1174]);
$fdisplay(file, "0x92E0,0x%h_0x%h", db_odd.mem_bank[1175],db_even.mem_bank[1175]);
$fdisplay(file, "0x9300,0x%h_0x%h", db_odd.mem_bank[1176],db_even.mem_bank[1176]);
$fdisplay(file, "0x9320,0x%h_0x%h", db_odd.mem_bank[1177],db_even.mem_bank[1177]);
$fdisplay(file, "0x9340,0x%h_0x%h", db_odd.mem_bank[1178],db_even.mem_bank[1178]);
$fdisplay(file, "0x9360,0x%h_0x%h", db_odd.mem_bank[1179],db_even.mem_bank[1179]);
$fdisplay(file, "0x9380,0x%h_0x%h", db_odd.mem_bank[1180],db_even.mem_bank[1180]);
$fdisplay(file, "0x93A0,0x%h_0x%h", db_odd.mem_bank[1181],db_even.mem_bank[1181]);
$fdisplay(file, "0x93C0,0x%h_0x%h", db_odd.mem_bank[1182],db_even.mem_bank[1182]);
$fdisplay(file, "0x93E0,0x%h_0x%h", db_odd.mem_bank[1183],db_even.mem_bank[1183]);
$fdisplay(file, "0x9400,0x%h_0x%h", db_odd.mem_bank[1184],db_even.mem_bank[1184]);
$fdisplay(file, "0x9420,0x%h_0x%h", db_odd.mem_bank[1185],db_even.mem_bank[1185]);
$fdisplay(file, "0x9440,0x%h_0x%h", db_odd.mem_bank[1186],db_even.mem_bank[1186]);
$fdisplay(file, "0x9460,0x%h_0x%h", db_odd.mem_bank[1187],db_even.mem_bank[1187]);
$fdisplay(file, "0x9480,0x%h_0x%h", db_odd.mem_bank[1188],db_even.mem_bank[1188]);
$fdisplay(file, "0x94A0,0x%h_0x%h", db_odd.mem_bank[1189],db_even.mem_bank[1189]);
$fdisplay(file, "0x94C0,0x%h_0x%h", db_odd.mem_bank[1190],db_even.mem_bank[1190]);
$fdisplay(file, "0x94E0,0x%h_0x%h", db_odd.mem_bank[1191],db_even.mem_bank[1191]);
$fdisplay(file, "0x9500,0x%h_0x%h", db_odd.mem_bank[1192],db_even.mem_bank[1192]);
$fdisplay(file, "0x9520,0x%h_0x%h", db_odd.mem_bank[1193],db_even.mem_bank[1193]);
$fdisplay(file, "0x9540,0x%h_0x%h", db_odd.mem_bank[1194],db_even.mem_bank[1194]);
$fdisplay(file, "0x9560,0x%h_0x%h", db_odd.mem_bank[1195],db_even.mem_bank[1195]);
$fdisplay(file, "0x9580,0x%h_0x%h", db_odd.mem_bank[1196],db_even.mem_bank[1196]);
$fdisplay(file, "0x95A0,0x%h_0x%h", db_odd.mem_bank[1197],db_even.mem_bank[1197]);
$fdisplay(file, "0x95C0,0x%h_0x%h", db_odd.mem_bank[1198],db_even.mem_bank[1198]);
$fdisplay(file, "0x95E0,0x%h_0x%h", db_odd.mem_bank[1199],db_even.mem_bank[1199]);
$fdisplay(file, "0x9600,0x%h_0x%h", db_odd.mem_bank[1200],db_even.mem_bank[1200]);
$fdisplay(file, "0x9620,0x%h_0x%h", db_odd.mem_bank[1201],db_even.mem_bank[1201]);
$fdisplay(file, "0x9640,0x%h_0x%h", db_odd.mem_bank[1202],db_even.mem_bank[1202]);
$fdisplay(file, "0x9660,0x%h_0x%h", db_odd.mem_bank[1203],db_even.mem_bank[1203]);
$fdisplay(file, "0x9680,0x%h_0x%h", db_odd.mem_bank[1204],db_even.mem_bank[1204]);
$fdisplay(file, "0x96A0,0x%h_0x%h", db_odd.mem_bank[1205],db_even.mem_bank[1205]);
$fdisplay(file, "0x96C0,0x%h_0x%h", db_odd.mem_bank[1206],db_even.mem_bank[1206]);
$fdisplay(file, "0x96E0,0x%h_0x%h", db_odd.mem_bank[1207],db_even.mem_bank[1207]);
$fdisplay(file, "0x9700,0x%h_0x%h", db_odd.mem_bank[1208],db_even.mem_bank[1208]);
$fdisplay(file, "0x9720,0x%h_0x%h", db_odd.mem_bank[1209],db_even.mem_bank[1209]);
$fdisplay(file, "0x9740,0x%h_0x%h", db_odd.mem_bank[1210],db_even.mem_bank[1210]);
$fdisplay(file, "0x9760,0x%h_0x%h", db_odd.mem_bank[1211],db_even.mem_bank[1211]);
$fdisplay(file, "0x9780,0x%h_0x%h", db_odd.mem_bank[1212],db_even.mem_bank[1212]);
$fdisplay(file, "0x97A0,0x%h_0x%h", db_odd.mem_bank[1213],db_even.mem_bank[1213]);
$fdisplay(file, "0x97C0,0x%h_0x%h", db_odd.mem_bank[1214],db_even.mem_bank[1214]);
$fdisplay(file, "0x97E0,0x%h_0x%h", db_odd.mem_bank[1215],db_even.mem_bank[1215]);
$fdisplay(file, "0x9800,0x%h_0x%h", db_odd.mem_bank[1216],db_even.mem_bank[1216]);
$fdisplay(file, "0x9820,0x%h_0x%h", db_odd.mem_bank[1217],db_even.mem_bank[1217]);
$fdisplay(file, "0x9840,0x%h_0x%h", db_odd.mem_bank[1218],db_even.mem_bank[1218]);
$fdisplay(file, "0x9860,0x%h_0x%h", db_odd.mem_bank[1219],db_even.mem_bank[1219]);
$fdisplay(file, "0x9880,0x%h_0x%h", db_odd.mem_bank[1220],db_even.mem_bank[1220]);
$fdisplay(file, "0x98A0,0x%h_0x%h", db_odd.mem_bank[1221],db_even.mem_bank[1221]);
$fdisplay(file, "0x98C0,0x%h_0x%h", db_odd.mem_bank[1222],db_even.mem_bank[1222]);
$fdisplay(file, "0x98E0,0x%h_0x%h", db_odd.mem_bank[1223],db_even.mem_bank[1223]);
$fdisplay(file, "0x9900,0x%h_0x%h", db_odd.mem_bank[1224],db_even.mem_bank[1224]);
$fdisplay(file, "0x9920,0x%h_0x%h", db_odd.mem_bank[1225],db_even.mem_bank[1225]);
$fdisplay(file, "0x9940,0x%h_0x%h", db_odd.mem_bank[1226],db_even.mem_bank[1226]);
$fdisplay(file, "0x9960,0x%h_0x%h", db_odd.mem_bank[1227],db_even.mem_bank[1227]);
$fdisplay(file, "0x9980,0x%h_0x%h", db_odd.mem_bank[1228],db_even.mem_bank[1228]);
$fdisplay(file, "0x99A0,0x%h_0x%h", db_odd.mem_bank[1229],db_even.mem_bank[1229]);
$fdisplay(file, "0x99C0,0x%h_0x%h", db_odd.mem_bank[1230],db_even.mem_bank[1230]);
$fdisplay(file, "0x99E0,0x%h_0x%h", db_odd.mem_bank[1231],db_even.mem_bank[1231]);
$fdisplay(file, "0x9A00,0x%h_0x%h", db_odd.mem_bank[1232],db_even.mem_bank[1232]);
$fdisplay(file, "0x9A20,0x%h_0x%h", db_odd.mem_bank[1233],db_even.mem_bank[1233]);
$fdisplay(file, "0x9A40,0x%h_0x%h", db_odd.mem_bank[1234],db_even.mem_bank[1234]);
$fdisplay(file, "0x9A60,0x%h_0x%h", db_odd.mem_bank[1235],db_even.mem_bank[1235]);
$fdisplay(file, "0x9A80,0x%h_0x%h", db_odd.mem_bank[1236],db_even.mem_bank[1236]);
$fdisplay(file, "0x9AA0,0x%h_0x%h", db_odd.mem_bank[1237],db_even.mem_bank[1237]);
$fdisplay(file, "0x9AC0,0x%h_0x%h", db_odd.mem_bank[1238],db_even.mem_bank[1238]);
$fdisplay(file, "0x9AE0,0x%h_0x%h", db_odd.mem_bank[1239],db_even.mem_bank[1239]);
$fdisplay(file, "0x9B00,0x%h_0x%h", db_odd.mem_bank[1240],db_even.mem_bank[1240]);
$fdisplay(file, "0x9B20,0x%h_0x%h", db_odd.mem_bank[1241],db_even.mem_bank[1241]);
$fdisplay(file, "0x9B40,0x%h_0x%h", db_odd.mem_bank[1242],db_even.mem_bank[1242]);
$fdisplay(file, "0x9B60,0x%h_0x%h", db_odd.mem_bank[1243],db_even.mem_bank[1243]);
$fdisplay(file, "0x9B80,0x%h_0x%h", db_odd.mem_bank[1244],db_even.mem_bank[1244]);
$fdisplay(file, "0x9BA0,0x%h_0x%h", db_odd.mem_bank[1245],db_even.mem_bank[1245]);
$fdisplay(file, "0x9BC0,0x%h_0x%h", db_odd.mem_bank[1246],db_even.mem_bank[1246]);
$fdisplay(file, "0x9BE0,0x%h_0x%h", db_odd.mem_bank[1247],db_even.mem_bank[1247]);
$fdisplay(file, "0x9C00,0x%h_0x%h", db_odd.mem_bank[1248],db_even.mem_bank[1248]);
$fdisplay(file, "0x9C20,0x%h_0x%h", db_odd.mem_bank[1249],db_even.mem_bank[1249]);
$fdisplay(file, "0x9C40,0x%h_0x%h", db_odd.mem_bank[1250],db_even.mem_bank[1250]);
$fdisplay(file, "0x9C60,0x%h_0x%h", db_odd.mem_bank[1251],db_even.mem_bank[1251]);
$fdisplay(file, "0x9C80,0x%h_0x%h", db_odd.mem_bank[1252],db_even.mem_bank[1252]);
$fdisplay(file, "0x9CA0,0x%h_0x%h", db_odd.mem_bank[1253],db_even.mem_bank[1253]);
$fdisplay(file, "0x9CC0,0x%h_0x%h", db_odd.mem_bank[1254],db_even.mem_bank[1254]);
$fdisplay(file, "0x9CE0,0x%h_0x%h", db_odd.mem_bank[1255],db_even.mem_bank[1255]);
$fdisplay(file, "0x9D00,0x%h_0x%h", db_odd.mem_bank[1256],db_even.mem_bank[1256]);
$fdisplay(file, "0x9D20,0x%h_0x%h", db_odd.mem_bank[1257],db_even.mem_bank[1257]);
$fdisplay(file, "0x9D40,0x%h_0x%h", db_odd.mem_bank[1258],db_even.mem_bank[1258]);
$fdisplay(file, "0x9D60,0x%h_0x%h", db_odd.mem_bank[1259],db_even.mem_bank[1259]);
$fdisplay(file, "0x9D80,0x%h_0x%h", db_odd.mem_bank[1260],db_even.mem_bank[1260]);
$fdisplay(file, "0x9DA0,0x%h_0x%h", db_odd.mem_bank[1261],db_even.mem_bank[1261]);
$fdisplay(file, "0x9DC0,0x%h_0x%h", db_odd.mem_bank[1262],db_even.mem_bank[1262]);
$fdisplay(file, "0x9DE0,0x%h_0x%h", db_odd.mem_bank[1263],db_even.mem_bank[1263]);
$fdisplay(file, "0x9E00,0x%h_0x%h", db_odd.mem_bank[1264],db_even.mem_bank[1264]);
$fdisplay(file, "0x9E20,0x%h_0x%h", db_odd.mem_bank[1265],db_even.mem_bank[1265]);
$fdisplay(file, "0x9E40,0x%h_0x%h", db_odd.mem_bank[1266],db_even.mem_bank[1266]);
$fdisplay(file, "0x9E60,0x%h_0x%h", db_odd.mem_bank[1267],db_even.mem_bank[1267]);
$fdisplay(file, "0x9E80,0x%h_0x%h", db_odd.mem_bank[1268],db_even.mem_bank[1268]);
$fdisplay(file, "0x9EA0,0x%h_0x%h", db_odd.mem_bank[1269],db_even.mem_bank[1269]);
$fdisplay(file, "0x9EC0,0x%h_0x%h", db_odd.mem_bank[1270],db_even.mem_bank[1270]);
$fdisplay(file, "0x9EE0,0x%h_0x%h", db_odd.mem_bank[1271],db_even.mem_bank[1271]);
$fdisplay(file, "0x9F00,0x%h_0x%h", db_odd.mem_bank[1272],db_even.mem_bank[1272]);
$fdisplay(file, "0x9F20,0x%h_0x%h", db_odd.mem_bank[1273],db_even.mem_bank[1273]);
$fdisplay(file, "0x9F40,0x%h_0x%h", db_odd.mem_bank[1274],db_even.mem_bank[1274]);
$fdisplay(file, "0x9F60,0x%h_0x%h", db_odd.mem_bank[1275],db_even.mem_bank[1275]);
$fdisplay(file, "0x9F80,0x%h_0x%h", db_odd.mem_bank[1276],db_even.mem_bank[1276]);
$fdisplay(file, "0x9FA0,0x%h_0x%h", db_odd.mem_bank[1277],db_even.mem_bank[1277]);
$fdisplay(file, "0x9FC0,0x%h_0x%h", db_odd.mem_bank[1278],db_even.mem_bank[1278]);
$fdisplay(file, "0x9FE0,0x%h_0x%h", db_odd.mem_bank[1279],db_even.mem_bank[1279]);
$fdisplay(file, "0xA000,0x%h_0x%h", db_odd.mem_bank[1280],db_even.mem_bank[1280]);
$fdisplay(file, "0xA020,0x%h_0x%h", db_odd.mem_bank[1281],db_even.mem_bank[1281]);
$fdisplay(file, "0xA040,0x%h_0x%h", db_odd.mem_bank[1282],db_even.mem_bank[1282]);
$fdisplay(file, "0xA060,0x%h_0x%h", db_odd.mem_bank[1283],db_even.mem_bank[1283]);
$fdisplay(file, "0xA080,0x%h_0x%h", db_odd.mem_bank[1284],db_even.mem_bank[1284]);
$fdisplay(file, "0xA0A0,0x%h_0x%h", db_odd.mem_bank[1285],db_even.mem_bank[1285]);
$fdisplay(file, "0xA0C0,0x%h_0x%h", db_odd.mem_bank[1286],db_even.mem_bank[1286]);
$fdisplay(file, "0xA0E0,0x%h_0x%h", db_odd.mem_bank[1287],db_even.mem_bank[1287]);
$fdisplay(file, "0xA100,0x%h_0x%h", db_odd.mem_bank[1288],db_even.mem_bank[1288]);
$fdisplay(file, "0xA120,0x%h_0x%h", db_odd.mem_bank[1289],db_even.mem_bank[1289]);
$fdisplay(file, "0xA140,0x%h_0x%h", db_odd.mem_bank[1290],db_even.mem_bank[1290]);
$fdisplay(file, "0xA160,0x%h_0x%h", db_odd.mem_bank[1291],db_even.mem_bank[1291]);
$fdisplay(file, "0xA180,0x%h_0x%h", db_odd.mem_bank[1292],db_even.mem_bank[1292]);
$fdisplay(file, "0xA1A0,0x%h_0x%h", db_odd.mem_bank[1293],db_even.mem_bank[1293]);
$fdisplay(file, "0xA1C0,0x%h_0x%h", db_odd.mem_bank[1294],db_even.mem_bank[1294]);
$fdisplay(file, "0xA1E0,0x%h_0x%h", db_odd.mem_bank[1295],db_even.mem_bank[1295]);
$fdisplay(file, "0xA200,0x%h_0x%h", db_odd.mem_bank[1296],db_even.mem_bank[1296]);
$fdisplay(file, "0xA220,0x%h_0x%h", db_odd.mem_bank[1297],db_even.mem_bank[1297]);
$fdisplay(file, "0xA240,0x%h_0x%h", db_odd.mem_bank[1298],db_even.mem_bank[1298]);
$fdisplay(file, "0xA260,0x%h_0x%h", db_odd.mem_bank[1299],db_even.mem_bank[1299]);
$fdisplay(file, "0xA280,0x%h_0x%h", db_odd.mem_bank[1300],db_even.mem_bank[1300]);
$fdisplay(file, "0xA2A0,0x%h_0x%h", db_odd.mem_bank[1301],db_even.mem_bank[1301]);
$fdisplay(file, "0xA2C0,0x%h_0x%h", db_odd.mem_bank[1302],db_even.mem_bank[1302]);
$fdisplay(file, "0xA2E0,0x%h_0x%h", db_odd.mem_bank[1303],db_even.mem_bank[1303]);
$fdisplay(file, "0xA300,0x%h_0x%h", db_odd.mem_bank[1304],db_even.mem_bank[1304]);
$fdisplay(file, "0xA320,0x%h_0x%h", db_odd.mem_bank[1305],db_even.mem_bank[1305]);
$fdisplay(file, "0xA340,0x%h_0x%h", db_odd.mem_bank[1306],db_even.mem_bank[1306]);
$fdisplay(file, "0xA360,0x%h_0x%h", db_odd.mem_bank[1307],db_even.mem_bank[1307]);
$fdisplay(file, "0xA380,0x%h_0x%h", db_odd.mem_bank[1308],db_even.mem_bank[1308]);
$fdisplay(file, "0xA3A0,0x%h_0x%h", db_odd.mem_bank[1309],db_even.mem_bank[1309]);
$fdisplay(file, "0xA3C0,0x%h_0x%h", db_odd.mem_bank[1310],db_even.mem_bank[1310]);
$fdisplay(file, "0xA3E0,0x%h_0x%h", db_odd.mem_bank[1311],db_even.mem_bank[1311]);
$fdisplay(file, "0xA400,0x%h_0x%h", db_odd.mem_bank[1312],db_even.mem_bank[1312]);
$fdisplay(file, "0xA420,0x%h_0x%h", db_odd.mem_bank[1313],db_even.mem_bank[1313]);
$fdisplay(file, "0xA440,0x%h_0x%h", db_odd.mem_bank[1314],db_even.mem_bank[1314]);
$fdisplay(file, "0xA460,0x%h_0x%h", db_odd.mem_bank[1315],db_even.mem_bank[1315]);
$fdisplay(file, "0xA480,0x%h_0x%h", db_odd.mem_bank[1316],db_even.mem_bank[1316]);
$fdisplay(file, "0xA4A0,0x%h_0x%h", db_odd.mem_bank[1317],db_even.mem_bank[1317]);
$fdisplay(file, "0xA4C0,0x%h_0x%h", db_odd.mem_bank[1318],db_even.mem_bank[1318]);
$fdisplay(file, "0xA4E0,0x%h_0x%h", db_odd.mem_bank[1319],db_even.mem_bank[1319]);
$fdisplay(file, "0xA500,0x%h_0x%h", db_odd.mem_bank[1320],db_even.mem_bank[1320]);
$fdisplay(file, "0xA520,0x%h_0x%h", db_odd.mem_bank[1321],db_even.mem_bank[1321]);
$fdisplay(file, "0xA540,0x%h_0x%h", db_odd.mem_bank[1322],db_even.mem_bank[1322]);
$fdisplay(file, "0xA560,0x%h_0x%h", db_odd.mem_bank[1323],db_even.mem_bank[1323]);
$fdisplay(file, "0xA580,0x%h_0x%h", db_odd.mem_bank[1324],db_even.mem_bank[1324]);
$fdisplay(file, "0xA5A0,0x%h_0x%h", db_odd.mem_bank[1325],db_even.mem_bank[1325]);
$fdisplay(file, "0xA5C0,0x%h_0x%h", db_odd.mem_bank[1326],db_even.mem_bank[1326]);
$fdisplay(file, "0xA5E0,0x%h_0x%h", db_odd.mem_bank[1327],db_even.mem_bank[1327]);
$fdisplay(file, "0xA600,0x%h_0x%h", db_odd.mem_bank[1328],db_even.mem_bank[1328]);
$fdisplay(file, "0xA620,0x%h_0x%h", db_odd.mem_bank[1329],db_even.mem_bank[1329]);
$fdisplay(file, "0xA640,0x%h_0x%h", db_odd.mem_bank[1330],db_even.mem_bank[1330]);
$fdisplay(file, "0xA660,0x%h_0x%h", db_odd.mem_bank[1331],db_even.mem_bank[1331]);
$fdisplay(file, "0xA680,0x%h_0x%h", db_odd.mem_bank[1332],db_even.mem_bank[1332]);
$fdisplay(file, "0xA6A0,0x%h_0x%h", db_odd.mem_bank[1333],db_even.mem_bank[1333]);
$fdisplay(file, "0xA6C0,0x%h_0x%h", db_odd.mem_bank[1334],db_even.mem_bank[1334]);
$fdisplay(file, "0xA6E0,0x%h_0x%h", db_odd.mem_bank[1335],db_even.mem_bank[1335]);
$fdisplay(file, "0xA700,0x%h_0x%h", db_odd.mem_bank[1336],db_even.mem_bank[1336]);
$fdisplay(file, "0xA720,0x%h_0x%h", db_odd.mem_bank[1337],db_even.mem_bank[1337]);
$fdisplay(file, "0xA740,0x%h_0x%h", db_odd.mem_bank[1338],db_even.mem_bank[1338]);
$fdisplay(file, "0xA760,0x%h_0x%h", db_odd.mem_bank[1339],db_even.mem_bank[1339]);
$fdisplay(file, "0xA780,0x%h_0x%h", db_odd.mem_bank[1340],db_even.mem_bank[1340]);
$fdisplay(file, "0xA7A0,0x%h_0x%h", db_odd.mem_bank[1341],db_even.mem_bank[1341]);
$fdisplay(file, "0xA7C0,0x%h_0x%h", db_odd.mem_bank[1342],db_even.mem_bank[1342]);
$fdisplay(file, "0xA7E0,0x%h_0x%h", db_odd.mem_bank[1343],db_even.mem_bank[1343]);
$fdisplay(file, "0xA800,0x%h_0x%h", db_odd.mem_bank[1344],db_even.mem_bank[1344]);
$fdisplay(file, "0xA820,0x%h_0x%h", db_odd.mem_bank[1345],db_even.mem_bank[1345]);
$fdisplay(file, "0xA840,0x%h_0x%h", db_odd.mem_bank[1346],db_even.mem_bank[1346]);
$fdisplay(file, "0xA860,0x%h_0x%h", db_odd.mem_bank[1347],db_even.mem_bank[1347]);
$fdisplay(file, "0xA880,0x%h_0x%h", db_odd.mem_bank[1348],db_even.mem_bank[1348]);
$fdisplay(file, "0xA8A0,0x%h_0x%h", db_odd.mem_bank[1349],db_even.mem_bank[1349]);
$fdisplay(file, "0xA8C0,0x%h_0x%h", db_odd.mem_bank[1350],db_even.mem_bank[1350]);
$fdisplay(file, "0xA8E0,0x%h_0x%h", db_odd.mem_bank[1351],db_even.mem_bank[1351]);
$fdisplay(file, "0xA900,0x%h_0x%h", db_odd.mem_bank[1352],db_even.mem_bank[1352]);
$fdisplay(file, "0xA920,0x%h_0x%h", db_odd.mem_bank[1353],db_even.mem_bank[1353]);
$fdisplay(file, "0xA940,0x%h_0x%h", db_odd.mem_bank[1354],db_even.mem_bank[1354]);
$fdisplay(file, "0xA960,0x%h_0x%h", db_odd.mem_bank[1355],db_even.mem_bank[1355]);
$fdisplay(file, "0xA980,0x%h_0x%h", db_odd.mem_bank[1356],db_even.mem_bank[1356]);
$fdisplay(file, "0xA9A0,0x%h_0x%h", db_odd.mem_bank[1357],db_even.mem_bank[1357]);
$fdisplay(file, "0xA9C0,0x%h_0x%h", db_odd.mem_bank[1358],db_even.mem_bank[1358]);
$fdisplay(file, "0xA9E0,0x%h_0x%h", db_odd.mem_bank[1359],db_even.mem_bank[1359]);
$fdisplay(file, "0xAA00,0x%h_0x%h", db_odd.mem_bank[1360],db_even.mem_bank[1360]);
$fdisplay(file, "0xAA20,0x%h_0x%h", db_odd.mem_bank[1361],db_even.mem_bank[1361]);
$fdisplay(file, "0xAA40,0x%h_0x%h", db_odd.mem_bank[1362],db_even.mem_bank[1362]);
$fdisplay(file, "0xAA60,0x%h_0x%h", db_odd.mem_bank[1363],db_even.mem_bank[1363]);
$fdisplay(file, "0xAA80,0x%h_0x%h", db_odd.mem_bank[1364],db_even.mem_bank[1364]);
$fdisplay(file, "0xAAA0,0x%h_0x%h", db_odd.mem_bank[1365],db_even.mem_bank[1365]);
$fdisplay(file, "0xAAC0,0x%h_0x%h", db_odd.mem_bank[1366],db_even.mem_bank[1366]);
$fdisplay(file, "0xAAE0,0x%h_0x%h", db_odd.mem_bank[1367],db_even.mem_bank[1367]);
$fdisplay(file, "0xAB00,0x%h_0x%h", db_odd.mem_bank[1368],db_even.mem_bank[1368]);
$fdisplay(file, "0xAB20,0x%h_0x%h", db_odd.mem_bank[1369],db_even.mem_bank[1369]);
$fdisplay(file, "0xAB40,0x%h_0x%h", db_odd.mem_bank[1370],db_even.mem_bank[1370]);
$fdisplay(file, "0xAB60,0x%h_0x%h", db_odd.mem_bank[1371],db_even.mem_bank[1371]);
$fdisplay(file, "0xAB80,0x%h_0x%h", db_odd.mem_bank[1372],db_even.mem_bank[1372]);
$fdisplay(file, "0xABA0,0x%h_0x%h", db_odd.mem_bank[1373],db_even.mem_bank[1373]);
$fdisplay(file, "0xABC0,0x%h_0x%h", db_odd.mem_bank[1374],db_even.mem_bank[1374]);
$fdisplay(file, "0xABE0,0x%h_0x%h", db_odd.mem_bank[1375],db_even.mem_bank[1375]);
$fdisplay(file, "0xAC00,0x%h_0x%h", db_odd.mem_bank[1376],db_even.mem_bank[1376]);
$fdisplay(file, "0xAC20,0x%h_0x%h", db_odd.mem_bank[1377],db_even.mem_bank[1377]);
$fdisplay(file, "0xAC40,0x%h_0x%h", db_odd.mem_bank[1378],db_even.mem_bank[1378]);
$fdisplay(file, "0xAC60,0x%h_0x%h", db_odd.mem_bank[1379],db_even.mem_bank[1379]);
$fdisplay(file, "0xAC80,0x%h_0x%h", db_odd.mem_bank[1380],db_even.mem_bank[1380]);
$fdisplay(file, "0xACA0,0x%h_0x%h", db_odd.mem_bank[1381],db_even.mem_bank[1381]);
$fdisplay(file, "0xACC0,0x%h_0x%h", db_odd.mem_bank[1382],db_even.mem_bank[1382]);
$fdisplay(file, "0xACE0,0x%h_0x%h", db_odd.mem_bank[1383],db_even.mem_bank[1383]);
$fdisplay(file, "0xAD00,0x%h_0x%h", db_odd.mem_bank[1384],db_even.mem_bank[1384]);
$fdisplay(file, "0xAD20,0x%h_0x%h", db_odd.mem_bank[1385],db_even.mem_bank[1385]);
$fdisplay(file, "0xAD40,0x%h_0x%h", db_odd.mem_bank[1386],db_even.mem_bank[1386]);
$fdisplay(file, "0xAD60,0x%h_0x%h", db_odd.mem_bank[1387],db_even.mem_bank[1387]);
$fdisplay(file, "0xAD80,0x%h_0x%h", db_odd.mem_bank[1388],db_even.mem_bank[1388]);
$fdisplay(file, "0xADA0,0x%h_0x%h", db_odd.mem_bank[1389],db_even.mem_bank[1389]);
$fdisplay(file, "0xADC0,0x%h_0x%h", db_odd.mem_bank[1390],db_even.mem_bank[1390]);
$fdisplay(file, "0xADE0,0x%h_0x%h", db_odd.mem_bank[1391],db_even.mem_bank[1391]);
$fdisplay(file, "0xAE00,0x%h_0x%h", db_odd.mem_bank[1392],db_even.mem_bank[1392]);
$fdisplay(file, "0xAE20,0x%h_0x%h", db_odd.mem_bank[1393],db_even.mem_bank[1393]);
$fdisplay(file, "0xAE40,0x%h_0x%h", db_odd.mem_bank[1394],db_even.mem_bank[1394]);
$fdisplay(file, "0xAE60,0x%h_0x%h", db_odd.mem_bank[1395],db_even.mem_bank[1395]);
$fdisplay(file, "0xAE80,0x%h_0x%h", db_odd.mem_bank[1396],db_even.mem_bank[1396]);
$fdisplay(file, "0xAEA0,0x%h_0x%h", db_odd.mem_bank[1397],db_even.mem_bank[1397]);
$fdisplay(file, "0xAEC0,0x%h_0x%h", db_odd.mem_bank[1398],db_even.mem_bank[1398]);
$fdisplay(file, "0xAEE0,0x%h_0x%h", db_odd.mem_bank[1399],db_even.mem_bank[1399]);
$fdisplay(file, "0xAF00,0x%h_0x%h", db_odd.mem_bank[1400],db_even.mem_bank[1400]);
$fdisplay(file, "0xAF20,0x%h_0x%h", db_odd.mem_bank[1401],db_even.mem_bank[1401]);
$fdisplay(file, "0xAF40,0x%h_0x%h", db_odd.mem_bank[1402],db_even.mem_bank[1402]);
$fdisplay(file, "0xAF60,0x%h_0x%h", db_odd.mem_bank[1403],db_even.mem_bank[1403]);
$fdisplay(file, "0xAF80,0x%h_0x%h", db_odd.mem_bank[1404],db_even.mem_bank[1404]);
$fdisplay(file, "0xAFA0,0x%h_0x%h", db_odd.mem_bank[1405],db_even.mem_bank[1405]);
$fdisplay(file, "0xAFC0,0x%h_0x%h", db_odd.mem_bank[1406],db_even.mem_bank[1406]);
$fdisplay(file, "0xAFE0,0x%h_0x%h", db_odd.mem_bank[1407],db_even.mem_bank[1407]);
$fdisplay(file, "0xB000,0x%h_0x%h", db_odd.mem_bank[1408],db_even.mem_bank[1408]);
$fdisplay(file, "0xB020,0x%h_0x%h", db_odd.mem_bank[1409],db_even.mem_bank[1409]);
$fdisplay(file, "0xB040,0x%h_0x%h", db_odd.mem_bank[1410],db_even.mem_bank[1410]);
$fdisplay(file, "0xB060,0x%h_0x%h", db_odd.mem_bank[1411],db_even.mem_bank[1411]);
$fdisplay(file, "0xB080,0x%h_0x%h", db_odd.mem_bank[1412],db_even.mem_bank[1412]);
$fdisplay(file, "0xB0A0,0x%h_0x%h", db_odd.mem_bank[1413],db_even.mem_bank[1413]);
$fdisplay(file, "0xB0C0,0x%h_0x%h", db_odd.mem_bank[1414],db_even.mem_bank[1414]);
$fdisplay(file, "0xB0E0,0x%h_0x%h", db_odd.mem_bank[1415],db_even.mem_bank[1415]);
$fdisplay(file, "0xB100,0x%h_0x%h", db_odd.mem_bank[1416],db_even.mem_bank[1416]);
$fdisplay(file, "0xB120,0x%h_0x%h", db_odd.mem_bank[1417],db_even.mem_bank[1417]);
$fdisplay(file, "0xB140,0x%h_0x%h", db_odd.mem_bank[1418],db_even.mem_bank[1418]);
$fdisplay(file, "0xB160,0x%h_0x%h", db_odd.mem_bank[1419],db_even.mem_bank[1419]);
$fdisplay(file, "0xB180,0x%h_0x%h", db_odd.mem_bank[1420],db_even.mem_bank[1420]);
$fdisplay(file, "0xB1A0,0x%h_0x%h", db_odd.mem_bank[1421],db_even.mem_bank[1421]);
$fdisplay(file, "0xB1C0,0x%h_0x%h", db_odd.mem_bank[1422],db_even.mem_bank[1422]);
$fdisplay(file, "0xB1E0,0x%h_0x%h", db_odd.mem_bank[1423],db_even.mem_bank[1423]);
$fdisplay(file, "0xB200,0x%h_0x%h", db_odd.mem_bank[1424],db_even.mem_bank[1424]);
$fdisplay(file, "0xB220,0x%h_0x%h", db_odd.mem_bank[1425],db_even.mem_bank[1425]);
$fdisplay(file, "0xB240,0x%h_0x%h", db_odd.mem_bank[1426],db_even.mem_bank[1426]);
$fdisplay(file, "0xB260,0x%h_0x%h", db_odd.mem_bank[1427],db_even.mem_bank[1427]);
$fdisplay(file, "0xB280,0x%h_0x%h", db_odd.mem_bank[1428],db_even.mem_bank[1428]);
$fdisplay(file, "0xB2A0,0x%h_0x%h", db_odd.mem_bank[1429],db_even.mem_bank[1429]);
$fdisplay(file, "0xB2C0,0x%h_0x%h", db_odd.mem_bank[1430],db_even.mem_bank[1430]);
$fdisplay(file, "0xB2E0,0x%h_0x%h", db_odd.mem_bank[1431],db_even.mem_bank[1431]);
$fdisplay(file, "0xB300,0x%h_0x%h", db_odd.mem_bank[1432],db_even.mem_bank[1432]);
$fdisplay(file, "0xB320,0x%h_0x%h", db_odd.mem_bank[1433],db_even.mem_bank[1433]);
$fdisplay(file, "0xB340,0x%h_0x%h", db_odd.mem_bank[1434],db_even.mem_bank[1434]);
$fdisplay(file, "0xB360,0x%h_0x%h", db_odd.mem_bank[1435],db_even.mem_bank[1435]);
$fdisplay(file, "0xB380,0x%h_0x%h", db_odd.mem_bank[1436],db_even.mem_bank[1436]);
$fdisplay(file, "0xB3A0,0x%h_0x%h", db_odd.mem_bank[1437],db_even.mem_bank[1437]);
$fdisplay(file, "0xB3C0,0x%h_0x%h", db_odd.mem_bank[1438],db_even.mem_bank[1438]);
$fdisplay(file, "0xB3E0,0x%h_0x%h", db_odd.mem_bank[1439],db_even.mem_bank[1439]);
$fdisplay(file, "0xB400,0x%h_0x%h", db_odd.mem_bank[1440],db_even.mem_bank[1440]);
$fdisplay(file, "0xB420,0x%h_0x%h", db_odd.mem_bank[1441],db_even.mem_bank[1441]);
$fdisplay(file, "0xB440,0x%h_0x%h", db_odd.mem_bank[1442],db_even.mem_bank[1442]);
$fdisplay(file, "0xB460,0x%h_0x%h", db_odd.mem_bank[1443],db_even.mem_bank[1443]);
$fdisplay(file, "0xB480,0x%h_0x%h", db_odd.mem_bank[1444],db_even.mem_bank[1444]);
$fdisplay(file, "0xB4A0,0x%h_0x%h", db_odd.mem_bank[1445],db_even.mem_bank[1445]);
$fdisplay(file, "0xB4C0,0x%h_0x%h", db_odd.mem_bank[1446],db_even.mem_bank[1446]);
$fdisplay(file, "0xB4E0,0x%h_0x%h", db_odd.mem_bank[1447],db_even.mem_bank[1447]);
$fdisplay(file, "0xB500,0x%h_0x%h", db_odd.mem_bank[1448],db_even.mem_bank[1448]);
$fdisplay(file, "0xB520,0x%h_0x%h", db_odd.mem_bank[1449],db_even.mem_bank[1449]);
$fdisplay(file, "0xB540,0x%h_0x%h", db_odd.mem_bank[1450],db_even.mem_bank[1450]);
$fdisplay(file, "0xB560,0x%h_0x%h", db_odd.mem_bank[1451],db_even.mem_bank[1451]);
$fdisplay(file, "0xB580,0x%h_0x%h", db_odd.mem_bank[1452],db_even.mem_bank[1452]);
$fdisplay(file, "0xB5A0,0x%h_0x%h", db_odd.mem_bank[1453],db_even.mem_bank[1453]);
$fdisplay(file, "0xB5C0,0x%h_0x%h", db_odd.mem_bank[1454],db_even.mem_bank[1454]);
$fdisplay(file, "0xB5E0,0x%h_0x%h", db_odd.mem_bank[1455],db_even.mem_bank[1455]);
$fdisplay(file, "0xB600,0x%h_0x%h", db_odd.mem_bank[1456],db_even.mem_bank[1456]);
$fdisplay(file, "0xB620,0x%h_0x%h", db_odd.mem_bank[1457],db_even.mem_bank[1457]);
$fdisplay(file, "0xB640,0x%h_0x%h", db_odd.mem_bank[1458],db_even.mem_bank[1458]);
$fdisplay(file, "0xB660,0x%h_0x%h", db_odd.mem_bank[1459],db_even.mem_bank[1459]);
$fdisplay(file, "0xB680,0x%h_0x%h", db_odd.mem_bank[1460],db_even.mem_bank[1460]);
$fdisplay(file, "0xB6A0,0x%h_0x%h", db_odd.mem_bank[1461],db_even.mem_bank[1461]);
$fdisplay(file, "0xB6C0,0x%h_0x%h", db_odd.mem_bank[1462],db_even.mem_bank[1462]);
$fdisplay(file, "0xB6E0,0x%h_0x%h", db_odd.mem_bank[1463],db_even.mem_bank[1463]);
$fdisplay(file, "0xB700,0x%h_0x%h", db_odd.mem_bank[1464],db_even.mem_bank[1464]);
$fdisplay(file, "0xB720,0x%h_0x%h", db_odd.mem_bank[1465],db_even.mem_bank[1465]);
$fdisplay(file, "0xB740,0x%h_0x%h", db_odd.mem_bank[1466],db_even.mem_bank[1466]);
$fdisplay(file, "0xB760,0x%h_0x%h", db_odd.mem_bank[1467],db_even.mem_bank[1467]);
$fdisplay(file, "0xB780,0x%h_0x%h", db_odd.mem_bank[1468],db_even.mem_bank[1468]);
$fdisplay(file, "0xB7A0,0x%h_0x%h", db_odd.mem_bank[1469],db_even.mem_bank[1469]);
$fdisplay(file, "0xB7C0,0x%h_0x%h", db_odd.mem_bank[1470],db_even.mem_bank[1470]);
$fdisplay(file, "0xB7E0,0x%h_0x%h", db_odd.mem_bank[1471],db_even.mem_bank[1471]);
$fdisplay(file, "0xB800,0x%h_0x%h", db_odd.mem_bank[1472],db_even.mem_bank[1472]);
$fdisplay(file, "0xB820,0x%h_0x%h", db_odd.mem_bank[1473],db_even.mem_bank[1473]);
$fdisplay(file, "0xB840,0x%h_0x%h", db_odd.mem_bank[1474],db_even.mem_bank[1474]);
$fdisplay(file, "0xB860,0x%h_0x%h", db_odd.mem_bank[1475],db_even.mem_bank[1475]);
$fdisplay(file, "0xB880,0x%h_0x%h", db_odd.mem_bank[1476],db_even.mem_bank[1476]);
$fdisplay(file, "0xB8A0,0x%h_0x%h", db_odd.mem_bank[1477],db_even.mem_bank[1477]);
$fdisplay(file, "0xB8C0,0x%h_0x%h", db_odd.mem_bank[1478],db_even.mem_bank[1478]);
$fdisplay(file, "0xB8E0,0x%h_0x%h", db_odd.mem_bank[1479],db_even.mem_bank[1479]);
$fdisplay(file, "0xB900,0x%h_0x%h", db_odd.mem_bank[1480],db_even.mem_bank[1480]);
$fdisplay(file, "0xB920,0x%h_0x%h", db_odd.mem_bank[1481],db_even.mem_bank[1481]);
$fdisplay(file, "0xB940,0x%h_0x%h", db_odd.mem_bank[1482],db_even.mem_bank[1482]);
$fdisplay(file, "0xB960,0x%h_0x%h", db_odd.mem_bank[1483],db_even.mem_bank[1483]);
$fdisplay(file, "0xB980,0x%h_0x%h", db_odd.mem_bank[1484],db_even.mem_bank[1484]);
$fdisplay(file, "0xB9A0,0x%h_0x%h", db_odd.mem_bank[1485],db_even.mem_bank[1485]);
$fdisplay(file, "0xB9C0,0x%h_0x%h", db_odd.mem_bank[1486],db_even.mem_bank[1486]);
$fdisplay(file, "0xB9E0,0x%h_0x%h", db_odd.mem_bank[1487],db_even.mem_bank[1487]);
$fdisplay(file, "0xBA00,0x%h_0x%h", db_odd.mem_bank[1488],db_even.mem_bank[1488]);
$fdisplay(file, "0xBA20,0x%h_0x%h", db_odd.mem_bank[1489],db_even.mem_bank[1489]);
$fdisplay(file, "0xBA40,0x%h_0x%h", db_odd.mem_bank[1490],db_even.mem_bank[1490]);
$fdisplay(file, "0xBA60,0x%h_0x%h", db_odd.mem_bank[1491],db_even.mem_bank[1491]);
$fdisplay(file, "0xBA80,0x%h_0x%h", db_odd.mem_bank[1492],db_even.mem_bank[1492]);
$fdisplay(file, "0xBAA0,0x%h_0x%h", db_odd.mem_bank[1493],db_even.mem_bank[1493]);
$fdisplay(file, "0xBAC0,0x%h_0x%h", db_odd.mem_bank[1494],db_even.mem_bank[1494]);
$fdisplay(file, "0xBAE0,0x%h_0x%h", db_odd.mem_bank[1495],db_even.mem_bank[1495]);
$fdisplay(file, "0xBB00,0x%h_0x%h", db_odd.mem_bank[1496],db_even.mem_bank[1496]);
$fdisplay(file, "0xBB20,0x%h_0x%h", db_odd.mem_bank[1497],db_even.mem_bank[1497]);
$fdisplay(file, "0xBB40,0x%h_0x%h", db_odd.mem_bank[1498],db_even.mem_bank[1498]);
$fdisplay(file, "0xBB60,0x%h_0x%h", db_odd.mem_bank[1499],db_even.mem_bank[1499]);
$fdisplay(file, "0xBB80,0x%h_0x%h", db_odd.mem_bank[1500],db_even.mem_bank[1500]);
$fdisplay(file, "0xBBA0,0x%h_0x%h", db_odd.mem_bank[1501],db_even.mem_bank[1501]);
$fdisplay(file, "0xBBC0,0x%h_0x%h", db_odd.mem_bank[1502],db_even.mem_bank[1502]);
$fdisplay(file, "0xBBE0,0x%h_0x%h", db_odd.mem_bank[1503],db_even.mem_bank[1503]);
$fdisplay(file, "0xBC00,0x%h_0x%h", db_odd.mem_bank[1504],db_even.mem_bank[1504]);
$fdisplay(file, "0xBC20,0x%h_0x%h", db_odd.mem_bank[1505],db_even.mem_bank[1505]);
$fdisplay(file, "0xBC40,0x%h_0x%h", db_odd.mem_bank[1506],db_even.mem_bank[1506]);
$fdisplay(file, "0xBC60,0x%h_0x%h", db_odd.mem_bank[1507],db_even.mem_bank[1507]);
$fdisplay(file, "0xBC80,0x%h_0x%h", db_odd.mem_bank[1508],db_even.mem_bank[1508]);
$fdisplay(file, "0xBCA0,0x%h_0x%h", db_odd.mem_bank[1509],db_even.mem_bank[1509]);
$fdisplay(file, "0xBCC0,0x%h_0x%h", db_odd.mem_bank[1510],db_even.mem_bank[1510]);
$fdisplay(file, "0xBCE0,0x%h_0x%h", db_odd.mem_bank[1511],db_even.mem_bank[1511]);
$fdisplay(file, "0xBD00,0x%h_0x%h", db_odd.mem_bank[1512],db_even.mem_bank[1512]);
$fdisplay(file, "0xBD20,0x%h_0x%h", db_odd.mem_bank[1513],db_even.mem_bank[1513]);
$fdisplay(file, "0xBD40,0x%h_0x%h", db_odd.mem_bank[1514],db_even.mem_bank[1514]);
$fdisplay(file, "0xBD60,0x%h_0x%h", db_odd.mem_bank[1515],db_even.mem_bank[1515]);
$fdisplay(file, "0xBD80,0x%h_0x%h", db_odd.mem_bank[1516],db_even.mem_bank[1516]);
$fdisplay(file, "0xBDA0,0x%h_0x%h", db_odd.mem_bank[1517],db_even.mem_bank[1517]);
$fdisplay(file, "0xBDC0,0x%h_0x%h", db_odd.mem_bank[1518],db_even.mem_bank[1518]);
$fdisplay(file, "0xBDE0,0x%h_0x%h", db_odd.mem_bank[1519],db_even.mem_bank[1519]);
$fdisplay(file, "0xBE00,0x%h_0x%h", db_odd.mem_bank[1520],db_even.mem_bank[1520]);
$fdisplay(file, "0xBE20,0x%h_0x%h", db_odd.mem_bank[1521],db_even.mem_bank[1521]);
$fdisplay(file, "0xBE40,0x%h_0x%h", db_odd.mem_bank[1522],db_even.mem_bank[1522]);
$fdisplay(file, "0xBE60,0x%h_0x%h", db_odd.mem_bank[1523],db_even.mem_bank[1523]);
$fdisplay(file, "0xBE80,0x%h_0x%h", db_odd.mem_bank[1524],db_even.mem_bank[1524]);
$fdisplay(file, "0xBEA0,0x%h_0x%h", db_odd.mem_bank[1525],db_even.mem_bank[1525]);
$fdisplay(file, "0xBEC0,0x%h_0x%h", db_odd.mem_bank[1526],db_even.mem_bank[1526]);
$fdisplay(file, "0xBEE0,0x%h_0x%h", db_odd.mem_bank[1527],db_even.mem_bank[1527]);
$fdisplay(file, "0xBF00,0x%h_0x%h", db_odd.mem_bank[1528],db_even.mem_bank[1528]);
$fdisplay(file, "0xBF20,0x%h_0x%h", db_odd.mem_bank[1529],db_even.mem_bank[1529]);
$fdisplay(file, "0xBF40,0x%h_0x%h", db_odd.mem_bank[1530],db_even.mem_bank[1530]);
$fdisplay(file, "0xBF60,0x%h_0x%h", db_odd.mem_bank[1531],db_even.mem_bank[1531]);
$fdisplay(file, "0xBF80,0x%h_0x%h", db_odd.mem_bank[1532],db_even.mem_bank[1532]);
$fdisplay(file, "0xBFA0,0x%h_0x%h", db_odd.mem_bank[1533],db_even.mem_bank[1533]);
$fdisplay(file, "0xBFC0,0x%h_0x%h", db_odd.mem_bank[1534],db_even.mem_bank[1534]);
$fdisplay(file, "0xBFE0,0x%h_0x%h", db_odd.mem_bank[1535],db_even.mem_bank[1535]);
$fdisplay(file, "0xC000,0x%h_0x%h", db_odd.mem_bank[1536],db_even.mem_bank[1536]);
$fdisplay(file, "0xC020,0x%h_0x%h", db_odd.mem_bank[1537],db_even.mem_bank[1537]);
$fdisplay(file, "0xC040,0x%h_0x%h", db_odd.mem_bank[1538],db_even.mem_bank[1538]);
$fdisplay(file, "0xC060,0x%h_0x%h", db_odd.mem_bank[1539],db_even.mem_bank[1539]);
$fdisplay(file, "0xC080,0x%h_0x%h", db_odd.mem_bank[1540],db_even.mem_bank[1540]);
$fdisplay(file, "0xC0A0,0x%h_0x%h", db_odd.mem_bank[1541],db_even.mem_bank[1541]);
$fdisplay(file, "0xC0C0,0x%h_0x%h", db_odd.mem_bank[1542],db_even.mem_bank[1542]);
$fdisplay(file, "0xC0E0,0x%h_0x%h", db_odd.mem_bank[1543],db_even.mem_bank[1543]);
$fdisplay(file, "0xC100,0x%h_0x%h", db_odd.mem_bank[1544],db_even.mem_bank[1544]);
$fdisplay(file, "0xC120,0x%h_0x%h", db_odd.mem_bank[1545],db_even.mem_bank[1545]);
$fdisplay(file, "0xC140,0x%h_0x%h", db_odd.mem_bank[1546],db_even.mem_bank[1546]);
$fdisplay(file, "0xC160,0x%h_0x%h", db_odd.mem_bank[1547],db_even.mem_bank[1547]);
$fdisplay(file, "0xC180,0x%h_0x%h", db_odd.mem_bank[1548],db_even.mem_bank[1548]);
$fdisplay(file, "0xC1A0,0x%h_0x%h", db_odd.mem_bank[1549],db_even.mem_bank[1549]);
$fdisplay(file, "0xC1C0,0x%h_0x%h", db_odd.mem_bank[1550],db_even.mem_bank[1550]);
$fdisplay(file, "0xC1E0,0x%h_0x%h", db_odd.mem_bank[1551],db_even.mem_bank[1551]);
$fdisplay(file, "0xC200,0x%h_0x%h", db_odd.mem_bank[1552],db_even.mem_bank[1552]);
$fdisplay(file, "0xC220,0x%h_0x%h", db_odd.mem_bank[1553],db_even.mem_bank[1553]);
$fdisplay(file, "0xC240,0x%h_0x%h", db_odd.mem_bank[1554],db_even.mem_bank[1554]);
$fdisplay(file, "0xC260,0x%h_0x%h", db_odd.mem_bank[1555],db_even.mem_bank[1555]);
$fdisplay(file, "0xC280,0x%h_0x%h", db_odd.mem_bank[1556],db_even.mem_bank[1556]);
$fdisplay(file, "0xC2A0,0x%h_0x%h", db_odd.mem_bank[1557],db_even.mem_bank[1557]);
$fdisplay(file, "0xC2C0,0x%h_0x%h", db_odd.mem_bank[1558],db_even.mem_bank[1558]);
$fdisplay(file, "0xC2E0,0x%h_0x%h", db_odd.mem_bank[1559],db_even.mem_bank[1559]);
$fdisplay(file, "0xC300,0x%h_0x%h", db_odd.mem_bank[1560],db_even.mem_bank[1560]);
$fdisplay(file, "0xC320,0x%h_0x%h", db_odd.mem_bank[1561],db_even.mem_bank[1561]);
$fdisplay(file, "0xC340,0x%h_0x%h", db_odd.mem_bank[1562],db_even.mem_bank[1562]);
$fdisplay(file, "0xC360,0x%h_0x%h", db_odd.mem_bank[1563],db_even.mem_bank[1563]);
$fdisplay(file, "0xC380,0x%h_0x%h", db_odd.mem_bank[1564],db_even.mem_bank[1564]);
$fdisplay(file, "0xC3A0,0x%h_0x%h", db_odd.mem_bank[1565],db_even.mem_bank[1565]);
$fdisplay(file, "0xC3C0,0x%h_0x%h", db_odd.mem_bank[1566],db_even.mem_bank[1566]);
$fdisplay(file, "0xC3E0,0x%h_0x%h", db_odd.mem_bank[1567],db_even.mem_bank[1567]);
$fdisplay(file, "0xC400,0x%h_0x%h", db_odd.mem_bank[1568],db_even.mem_bank[1568]);
$fdisplay(file, "0xC420,0x%h_0x%h", db_odd.mem_bank[1569],db_even.mem_bank[1569]);
$fdisplay(file, "0xC440,0x%h_0x%h", db_odd.mem_bank[1570],db_even.mem_bank[1570]);
$fdisplay(file, "0xC460,0x%h_0x%h", db_odd.mem_bank[1571],db_even.mem_bank[1571]);
$fdisplay(file, "0xC480,0x%h_0x%h", db_odd.mem_bank[1572],db_even.mem_bank[1572]);
$fdisplay(file, "0xC4A0,0x%h_0x%h", db_odd.mem_bank[1573],db_even.mem_bank[1573]);
$fdisplay(file, "0xC4C0,0x%h_0x%h", db_odd.mem_bank[1574],db_even.mem_bank[1574]);
$fdisplay(file, "0xC4E0,0x%h_0x%h", db_odd.mem_bank[1575],db_even.mem_bank[1575]);
$fdisplay(file, "0xC500,0x%h_0x%h", db_odd.mem_bank[1576],db_even.mem_bank[1576]);
$fdisplay(file, "0xC520,0x%h_0x%h", db_odd.mem_bank[1577],db_even.mem_bank[1577]);
$fdisplay(file, "0xC540,0x%h_0x%h", db_odd.mem_bank[1578],db_even.mem_bank[1578]);
$fdisplay(file, "0xC560,0x%h_0x%h", db_odd.mem_bank[1579],db_even.mem_bank[1579]);
$fdisplay(file, "0xC580,0x%h_0x%h", db_odd.mem_bank[1580],db_even.mem_bank[1580]);
$fdisplay(file, "0xC5A0,0x%h_0x%h", db_odd.mem_bank[1581],db_even.mem_bank[1581]);
$fdisplay(file, "0xC5C0,0x%h_0x%h", db_odd.mem_bank[1582],db_even.mem_bank[1582]);
$fdisplay(file, "0xC5E0,0x%h_0x%h", db_odd.mem_bank[1583],db_even.mem_bank[1583]);
$fdisplay(file, "0xC600,0x%h_0x%h", db_odd.mem_bank[1584],db_even.mem_bank[1584]);
$fdisplay(file, "0xC620,0x%h_0x%h", db_odd.mem_bank[1585],db_even.mem_bank[1585]);
$fdisplay(file, "0xC640,0x%h_0x%h", db_odd.mem_bank[1586],db_even.mem_bank[1586]);
$fdisplay(file, "0xC660,0x%h_0x%h", db_odd.mem_bank[1587],db_even.mem_bank[1587]);
$fdisplay(file, "0xC680,0x%h_0x%h", db_odd.mem_bank[1588],db_even.mem_bank[1588]);
$fdisplay(file, "0xC6A0,0x%h_0x%h", db_odd.mem_bank[1589],db_even.mem_bank[1589]);
$fdisplay(file, "0xC6C0,0x%h_0x%h", db_odd.mem_bank[1590],db_even.mem_bank[1590]);
$fdisplay(file, "0xC6E0,0x%h_0x%h", db_odd.mem_bank[1591],db_even.mem_bank[1591]);
$fdisplay(file, "0xC700,0x%h_0x%h", db_odd.mem_bank[1592],db_even.mem_bank[1592]);
$fdisplay(file, "0xC720,0x%h_0x%h", db_odd.mem_bank[1593],db_even.mem_bank[1593]);
$fdisplay(file, "0xC740,0x%h_0x%h", db_odd.mem_bank[1594],db_even.mem_bank[1594]);
$fdisplay(file, "0xC760,0x%h_0x%h", db_odd.mem_bank[1595],db_even.mem_bank[1595]);
$fdisplay(file, "0xC780,0x%h_0x%h", db_odd.mem_bank[1596],db_even.mem_bank[1596]);
$fdisplay(file, "0xC7A0,0x%h_0x%h", db_odd.mem_bank[1597],db_even.mem_bank[1597]);
$fdisplay(file, "0xC7C0,0x%h_0x%h", db_odd.mem_bank[1598],db_even.mem_bank[1598]);
$fdisplay(file, "0xC7E0,0x%h_0x%h", db_odd.mem_bank[1599],db_even.mem_bank[1599]);
$fdisplay(file, "0xC800,0x%h_0x%h", db_odd.mem_bank[1600],db_even.mem_bank[1600]);
$fdisplay(file, "0xC820,0x%h_0x%h", db_odd.mem_bank[1601],db_even.mem_bank[1601]);
$fdisplay(file, "0xC840,0x%h_0x%h", db_odd.mem_bank[1602],db_even.mem_bank[1602]);
$fdisplay(file, "0xC860,0x%h_0x%h", db_odd.mem_bank[1603],db_even.mem_bank[1603]);
$fdisplay(file, "0xC880,0x%h_0x%h", db_odd.mem_bank[1604],db_even.mem_bank[1604]);
$fdisplay(file, "0xC8A0,0x%h_0x%h", db_odd.mem_bank[1605],db_even.mem_bank[1605]);
$fdisplay(file, "0xC8C0,0x%h_0x%h", db_odd.mem_bank[1606],db_even.mem_bank[1606]);
$fdisplay(file, "0xC8E0,0x%h_0x%h", db_odd.mem_bank[1607],db_even.mem_bank[1607]);
$fdisplay(file, "0xC900,0x%h_0x%h", db_odd.mem_bank[1608],db_even.mem_bank[1608]);
$fdisplay(file, "0xC920,0x%h_0x%h", db_odd.mem_bank[1609],db_even.mem_bank[1609]);
$fdisplay(file, "0xC940,0x%h_0x%h", db_odd.mem_bank[1610],db_even.mem_bank[1610]);
$fdisplay(file, "0xC960,0x%h_0x%h", db_odd.mem_bank[1611],db_even.mem_bank[1611]);
$fdisplay(file, "0xC980,0x%h_0x%h", db_odd.mem_bank[1612],db_even.mem_bank[1612]);
$fdisplay(file, "0xC9A0,0x%h_0x%h", db_odd.mem_bank[1613],db_even.mem_bank[1613]);
$fdisplay(file, "0xC9C0,0x%h_0x%h", db_odd.mem_bank[1614],db_even.mem_bank[1614]);
$fdisplay(file, "0xC9E0,0x%h_0x%h", db_odd.mem_bank[1615],db_even.mem_bank[1615]);
$fdisplay(file, "0xCA00,0x%h_0x%h", db_odd.mem_bank[1616],db_even.mem_bank[1616]);
$fdisplay(file, "0xCA20,0x%h_0x%h", db_odd.mem_bank[1617],db_even.mem_bank[1617]);
$fdisplay(file, "0xCA40,0x%h_0x%h", db_odd.mem_bank[1618],db_even.mem_bank[1618]);
$fdisplay(file, "0xCA60,0x%h_0x%h", db_odd.mem_bank[1619],db_even.mem_bank[1619]);
$fdisplay(file, "0xCA80,0x%h_0x%h", db_odd.mem_bank[1620],db_even.mem_bank[1620]);
$fdisplay(file, "0xCAA0,0x%h_0x%h", db_odd.mem_bank[1621],db_even.mem_bank[1621]);
$fdisplay(file, "0xCAC0,0x%h_0x%h", db_odd.mem_bank[1622],db_even.mem_bank[1622]);
$fdisplay(file, "0xCAE0,0x%h_0x%h", db_odd.mem_bank[1623],db_even.mem_bank[1623]);
$fdisplay(file, "0xCB00,0x%h_0x%h", db_odd.mem_bank[1624],db_even.mem_bank[1624]);
$fdisplay(file, "0xCB20,0x%h_0x%h", db_odd.mem_bank[1625],db_even.mem_bank[1625]);
$fdisplay(file, "0xCB40,0x%h_0x%h", db_odd.mem_bank[1626],db_even.mem_bank[1626]);
$fdisplay(file, "0xCB60,0x%h_0x%h", db_odd.mem_bank[1627],db_even.mem_bank[1627]);
$fdisplay(file, "0xCB80,0x%h_0x%h", db_odd.mem_bank[1628],db_even.mem_bank[1628]);
$fdisplay(file, "0xCBA0,0x%h_0x%h", db_odd.mem_bank[1629],db_even.mem_bank[1629]);
$fdisplay(file, "0xCBC0,0x%h_0x%h", db_odd.mem_bank[1630],db_even.mem_bank[1630]);
$fdisplay(file, "0xCBE0,0x%h_0x%h", db_odd.mem_bank[1631],db_even.mem_bank[1631]);
$fdisplay(file, "0xCC00,0x%h_0x%h", db_odd.mem_bank[1632],db_even.mem_bank[1632]);
$fdisplay(file, "0xCC20,0x%h_0x%h", db_odd.mem_bank[1633],db_even.mem_bank[1633]);
$fdisplay(file, "0xCC40,0x%h_0x%h", db_odd.mem_bank[1634],db_even.mem_bank[1634]);
$fdisplay(file, "0xCC60,0x%h_0x%h", db_odd.mem_bank[1635],db_even.mem_bank[1635]);
$fdisplay(file, "0xCC80,0x%h_0x%h", db_odd.mem_bank[1636],db_even.mem_bank[1636]);
$fdisplay(file, "0xCCA0,0x%h_0x%h", db_odd.mem_bank[1637],db_even.mem_bank[1637]);
$fdisplay(file, "0xCCC0,0x%h_0x%h", db_odd.mem_bank[1638],db_even.mem_bank[1638]);
$fdisplay(file, "0xCCE0,0x%h_0x%h", db_odd.mem_bank[1639],db_even.mem_bank[1639]);
$fdisplay(file, "0xCD00,0x%h_0x%h", db_odd.mem_bank[1640],db_even.mem_bank[1640]);
$fdisplay(file, "0xCD20,0x%h_0x%h", db_odd.mem_bank[1641],db_even.mem_bank[1641]);
$fdisplay(file, "0xCD40,0x%h_0x%h", db_odd.mem_bank[1642],db_even.mem_bank[1642]);
$fdisplay(file, "0xCD60,0x%h_0x%h", db_odd.mem_bank[1643],db_even.mem_bank[1643]);
$fdisplay(file, "0xCD80,0x%h_0x%h", db_odd.mem_bank[1644],db_even.mem_bank[1644]);
$fdisplay(file, "0xCDA0,0x%h_0x%h", db_odd.mem_bank[1645],db_even.mem_bank[1645]);
$fdisplay(file, "0xCDC0,0x%h_0x%h", db_odd.mem_bank[1646],db_even.mem_bank[1646]);
$fdisplay(file, "0xCDE0,0x%h_0x%h", db_odd.mem_bank[1647],db_even.mem_bank[1647]);
$fdisplay(file, "0xCE00,0x%h_0x%h", db_odd.mem_bank[1648],db_even.mem_bank[1648]);
$fdisplay(file, "0xCE20,0x%h_0x%h", db_odd.mem_bank[1649],db_even.mem_bank[1649]);
$fdisplay(file, "0xCE40,0x%h_0x%h", db_odd.mem_bank[1650],db_even.mem_bank[1650]);
$fdisplay(file, "0xCE60,0x%h_0x%h", db_odd.mem_bank[1651],db_even.mem_bank[1651]);
$fdisplay(file, "0xCE80,0x%h_0x%h", db_odd.mem_bank[1652],db_even.mem_bank[1652]);
$fdisplay(file, "0xCEA0,0x%h_0x%h", db_odd.mem_bank[1653],db_even.mem_bank[1653]);
$fdisplay(file, "0xCEC0,0x%h_0x%h", db_odd.mem_bank[1654],db_even.mem_bank[1654]);
$fdisplay(file, "0xCEE0,0x%h_0x%h", db_odd.mem_bank[1655],db_even.mem_bank[1655]);
$fdisplay(file, "0xCF00,0x%h_0x%h", db_odd.mem_bank[1656],db_even.mem_bank[1656]);
$fdisplay(file, "0xCF20,0x%h_0x%h", db_odd.mem_bank[1657],db_even.mem_bank[1657]);
$fdisplay(file, "0xCF40,0x%h_0x%h", db_odd.mem_bank[1658],db_even.mem_bank[1658]);
$fdisplay(file, "0xCF60,0x%h_0x%h", db_odd.mem_bank[1659],db_even.mem_bank[1659]);
$fdisplay(file, "0xCF80,0x%h_0x%h", db_odd.mem_bank[1660],db_even.mem_bank[1660]);
$fdisplay(file, "0xCFA0,0x%h_0x%h", db_odd.mem_bank[1661],db_even.mem_bank[1661]);
$fdisplay(file, "0xCFC0,0x%h_0x%h", db_odd.mem_bank[1662],db_even.mem_bank[1662]);
$fdisplay(file, "0xCFE0,0x%h_0x%h", db_odd.mem_bank[1663],db_even.mem_bank[1663]);
$fdisplay(file, "0xD000,0x%h_0x%h", db_odd.mem_bank[1664],db_even.mem_bank[1664]);
$fdisplay(file, "0xD020,0x%h_0x%h", db_odd.mem_bank[1665],db_even.mem_bank[1665]);
$fdisplay(file, "0xD040,0x%h_0x%h", db_odd.mem_bank[1666],db_even.mem_bank[1666]);
$fdisplay(file, "0xD060,0x%h_0x%h", db_odd.mem_bank[1667],db_even.mem_bank[1667]);
$fdisplay(file, "0xD080,0x%h_0x%h", db_odd.mem_bank[1668],db_even.mem_bank[1668]);
$fdisplay(file, "0xD0A0,0x%h_0x%h", db_odd.mem_bank[1669],db_even.mem_bank[1669]);
$fdisplay(file, "0xD0C0,0x%h_0x%h", db_odd.mem_bank[1670],db_even.mem_bank[1670]);
$fdisplay(file, "0xD0E0,0x%h_0x%h", db_odd.mem_bank[1671],db_even.mem_bank[1671]);
$fdisplay(file, "0xD100,0x%h_0x%h", db_odd.mem_bank[1672],db_even.mem_bank[1672]);
$fdisplay(file, "0xD120,0x%h_0x%h", db_odd.mem_bank[1673],db_even.mem_bank[1673]);
$fdisplay(file, "0xD140,0x%h_0x%h", db_odd.mem_bank[1674],db_even.mem_bank[1674]);
$fdisplay(file, "0xD160,0x%h_0x%h", db_odd.mem_bank[1675],db_even.mem_bank[1675]);
$fdisplay(file, "0xD180,0x%h_0x%h", db_odd.mem_bank[1676],db_even.mem_bank[1676]);
$fdisplay(file, "0xD1A0,0x%h_0x%h", db_odd.mem_bank[1677],db_even.mem_bank[1677]);
$fdisplay(file, "0xD1C0,0x%h_0x%h", db_odd.mem_bank[1678],db_even.mem_bank[1678]);
$fdisplay(file, "0xD1E0,0x%h_0x%h", db_odd.mem_bank[1679],db_even.mem_bank[1679]);
$fdisplay(file, "0xD200,0x%h_0x%h", db_odd.mem_bank[1680],db_even.mem_bank[1680]);
$fdisplay(file, "0xD220,0x%h_0x%h", db_odd.mem_bank[1681],db_even.mem_bank[1681]);
$fdisplay(file, "0xD240,0x%h_0x%h", db_odd.mem_bank[1682],db_even.mem_bank[1682]);
$fdisplay(file, "0xD260,0x%h_0x%h", db_odd.mem_bank[1683],db_even.mem_bank[1683]);
$fdisplay(file, "0xD280,0x%h_0x%h", db_odd.mem_bank[1684],db_even.mem_bank[1684]);
$fdisplay(file, "0xD2A0,0x%h_0x%h", db_odd.mem_bank[1685],db_even.mem_bank[1685]);
$fdisplay(file, "0xD2C0,0x%h_0x%h", db_odd.mem_bank[1686],db_even.mem_bank[1686]);
$fdisplay(file, "0xD2E0,0x%h_0x%h", db_odd.mem_bank[1687],db_even.mem_bank[1687]);
$fdisplay(file, "0xD300,0x%h_0x%h", db_odd.mem_bank[1688],db_even.mem_bank[1688]);
$fdisplay(file, "0xD320,0x%h_0x%h", db_odd.mem_bank[1689],db_even.mem_bank[1689]);
$fdisplay(file, "0xD340,0x%h_0x%h", db_odd.mem_bank[1690],db_even.mem_bank[1690]);
$fdisplay(file, "0xD360,0x%h_0x%h", db_odd.mem_bank[1691],db_even.mem_bank[1691]);
$fdisplay(file, "0xD380,0x%h_0x%h", db_odd.mem_bank[1692],db_even.mem_bank[1692]);
$fdisplay(file, "0xD3A0,0x%h_0x%h", db_odd.mem_bank[1693],db_even.mem_bank[1693]);
$fdisplay(file, "0xD3C0,0x%h_0x%h", db_odd.mem_bank[1694],db_even.mem_bank[1694]);
$fdisplay(file, "0xD3E0,0x%h_0x%h", db_odd.mem_bank[1695],db_even.mem_bank[1695]);
$fdisplay(file, "0xD400,0x%h_0x%h", db_odd.mem_bank[1696],db_even.mem_bank[1696]);
$fdisplay(file, "0xD420,0x%h_0x%h", db_odd.mem_bank[1697],db_even.mem_bank[1697]);
$fdisplay(file, "0xD440,0x%h_0x%h", db_odd.mem_bank[1698],db_even.mem_bank[1698]);
$fdisplay(file, "0xD460,0x%h_0x%h", db_odd.mem_bank[1699],db_even.mem_bank[1699]);
$fdisplay(file, "0xD480,0x%h_0x%h", db_odd.mem_bank[1700],db_even.mem_bank[1700]);
$fdisplay(file, "0xD4A0,0x%h_0x%h", db_odd.mem_bank[1701],db_even.mem_bank[1701]);
$fdisplay(file, "0xD4C0,0x%h_0x%h", db_odd.mem_bank[1702],db_even.mem_bank[1702]);
$fdisplay(file, "0xD4E0,0x%h_0x%h", db_odd.mem_bank[1703],db_even.mem_bank[1703]);
$fdisplay(file, "0xD500,0x%h_0x%h", db_odd.mem_bank[1704],db_even.mem_bank[1704]);
$fdisplay(file, "0xD520,0x%h_0x%h", db_odd.mem_bank[1705],db_even.mem_bank[1705]);
$fdisplay(file, "0xD540,0x%h_0x%h", db_odd.mem_bank[1706],db_even.mem_bank[1706]);
$fdisplay(file, "0xD560,0x%h_0x%h", db_odd.mem_bank[1707],db_even.mem_bank[1707]);
$fdisplay(file, "0xD580,0x%h_0x%h", db_odd.mem_bank[1708],db_even.mem_bank[1708]);
$fdisplay(file, "0xD5A0,0x%h_0x%h", db_odd.mem_bank[1709],db_even.mem_bank[1709]);
$fdisplay(file, "0xD5C0,0x%h_0x%h", db_odd.mem_bank[1710],db_even.mem_bank[1710]);
$fdisplay(file, "0xD5E0,0x%h_0x%h", db_odd.mem_bank[1711],db_even.mem_bank[1711]);
$fdisplay(file, "0xD600,0x%h_0x%h", db_odd.mem_bank[1712],db_even.mem_bank[1712]);
$fdisplay(file, "0xD620,0x%h_0x%h", db_odd.mem_bank[1713],db_even.mem_bank[1713]);
$fdisplay(file, "0xD640,0x%h_0x%h", db_odd.mem_bank[1714],db_even.mem_bank[1714]);
$fdisplay(file, "0xD660,0x%h_0x%h", db_odd.mem_bank[1715],db_even.mem_bank[1715]);
$fdisplay(file, "0xD680,0x%h_0x%h", db_odd.mem_bank[1716],db_even.mem_bank[1716]);
$fdisplay(file, "0xD6A0,0x%h_0x%h", db_odd.mem_bank[1717],db_even.mem_bank[1717]);
$fdisplay(file, "0xD6C0,0x%h_0x%h", db_odd.mem_bank[1718],db_even.mem_bank[1718]);
$fdisplay(file, "0xD6E0,0x%h_0x%h", db_odd.mem_bank[1719],db_even.mem_bank[1719]);
$fdisplay(file, "0xD700,0x%h_0x%h", db_odd.mem_bank[1720],db_even.mem_bank[1720]);
$fdisplay(file, "0xD720,0x%h_0x%h", db_odd.mem_bank[1721],db_even.mem_bank[1721]);
$fdisplay(file, "0xD740,0x%h_0x%h", db_odd.mem_bank[1722],db_even.mem_bank[1722]);
$fdisplay(file, "0xD760,0x%h_0x%h", db_odd.mem_bank[1723],db_even.mem_bank[1723]);
$fdisplay(file, "0xD780,0x%h_0x%h", db_odd.mem_bank[1724],db_even.mem_bank[1724]);
$fdisplay(file, "0xD7A0,0x%h_0x%h", db_odd.mem_bank[1725],db_even.mem_bank[1725]);
$fdisplay(file, "0xD7C0,0x%h_0x%h", db_odd.mem_bank[1726],db_even.mem_bank[1726]);
$fdisplay(file, "0xD7E0,0x%h_0x%h", db_odd.mem_bank[1727],db_even.mem_bank[1727]);
$fdisplay(file, "0xD800,0x%h_0x%h", db_odd.mem_bank[1728],db_even.mem_bank[1728]);
$fdisplay(file, "0xD820,0x%h_0x%h", db_odd.mem_bank[1729],db_even.mem_bank[1729]);
$fdisplay(file, "0xD840,0x%h_0x%h", db_odd.mem_bank[1730],db_even.mem_bank[1730]);
$fdisplay(file, "0xD860,0x%h_0x%h", db_odd.mem_bank[1731],db_even.mem_bank[1731]);
$fdisplay(file, "0xD880,0x%h_0x%h", db_odd.mem_bank[1732],db_even.mem_bank[1732]);
$fdisplay(file, "0xD8A0,0x%h_0x%h", db_odd.mem_bank[1733],db_even.mem_bank[1733]);
$fdisplay(file, "0xD8C0,0x%h_0x%h", db_odd.mem_bank[1734],db_even.mem_bank[1734]);
$fdisplay(file, "0xD8E0,0x%h_0x%h", db_odd.mem_bank[1735],db_even.mem_bank[1735]);
$fdisplay(file, "0xD900,0x%h_0x%h", db_odd.mem_bank[1736],db_even.mem_bank[1736]);
$fdisplay(file, "0xD920,0x%h_0x%h", db_odd.mem_bank[1737],db_even.mem_bank[1737]);
$fdisplay(file, "0xD940,0x%h_0x%h", db_odd.mem_bank[1738],db_even.mem_bank[1738]);
$fdisplay(file, "0xD960,0x%h_0x%h", db_odd.mem_bank[1739],db_even.mem_bank[1739]);
$fdisplay(file, "0xD980,0x%h_0x%h", db_odd.mem_bank[1740],db_even.mem_bank[1740]);
$fdisplay(file, "0xD9A0,0x%h_0x%h", db_odd.mem_bank[1741],db_even.mem_bank[1741]);
$fdisplay(file, "0xD9C0,0x%h_0x%h", db_odd.mem_bank[1742],db_even.mem_bank[1742]);
$fdisplay(file, "0xD9E0,0x%h_0x%h", db_odd.mem_bank[1743],db_even.mem_bank[1743]);
$fdisplay(file, "0xDA00,0x%h_0x%h", db_odd.mem_bank[1744],db_even.mem_bank[1744]);
$fdisplay(file, "0xDA20,0x%h_0x%h", db_odd.mem_bank[1745],db_even.mem_bank[1745]);
$fdisplay(file, "0xDA40,0x%h_0x%h", db_odd.mem_bank[1746],db_even.mem_bank[1746]);
$fdisplay(file, "0xDA60,0x%h_0x%h", db_odd.mem_bank[1747],db_even.mem_bank[1747]);
$fdisplay(file, "0xDA80,0x%h_0x%h", db_odd.mem_bank[1748],db_even.mem_bank[1748]);
$fdisplay(file, "0xDAA0,0x%h_0x%h", db_odd.mem_bank[1749],db_even.mem_bank[1749]);
$fdisplay(file, "0xDAC0,0x%h_0x%h", db_odd.mem_bank[1750],db_even.mem_bank[1750]);
$fdisplay(file, "0xDAE0,0x%h_0x%h", db_odd.mem_bank[1751],db_even.mem_bank[1751]);
$fdisplay(file, "0xDB00,0x%h_0x%h", db_odd.mem_bank[1752],db_even.mem_bank[1752]);
$fdisplay(file, "0xDB20,0x%h_0x%h", db_odd.mem_bank[1753],db_even.mem_bank[1753]);
$fdisplay(file, "0xDB40,0x%h_0x%h", db_odd.mem_bank[1754],db_even.mem_bank[1754]);
$fdisplay(file, "0xDB60,0x%h_0x%h", db_odd.mem_bank[1755],db_even.mem_bank[1755]);
$fdisplay(file, "0xDB80,0x%h_0x%h", db_odd.mem_bank[1756],db_even.mem_bank[1756]);
$fdisplay(file, "0xDBA0,0x%h_0x%h", db_odd.mem_bank[1757],db_even.mem_bank[1757]);
$fdisplay(file, "0xDBC0,0x%h_0x%h", db_odd.mem_bank[1758],db_even.mem_bank[1758]);
$fdisplay(file, "0xDBE0,0x%h_0x%h", db_odd.mem_bank[1759],db_even.mem_bank[1759]);
$fdisplay(file, "0xDC00,0x%h_0x%h", db_odd.mem_bank[1760],db_even.mem_bank[1760]);
$fdisplay(file, "0xDC20,0x%h_0x%h", db_odd.mem_bank[1761],db_even.mem_bank[1761]);
$fdisplay(file, "0xDC40,0x%h_0x%h", db_odd.mem_bank[1762],db_even.mem_bank[1762]);
$fdisplay(file, "0xDC60,0x%h_0x%h", db_odd.mem_bank[1763],db_even.mem_bank[1763]);
$fdisplay(file, "0xDC80,0x%h_0x%h", db_odd.mem_bank[1764],db_even.mem_bank[1764]);
$fdisplay(file, "0xDCA0,0x%h_0x%h", db_odd.mem_bank[1765],db_even.mem_bank[1765]);
$fdisplay(file, "0xDCC0,0x%h_0x%h", db_odd.mem_bank[1766],db_even.mem_bank[1766]);
$fdisplay(file, "0xDCE0,0x%h_0x%h", db_odd.mem_bank[1767],db_even.mem_bank[1767]);
$fdisplay(file, "0xDD00,0x%h_0x%h", db_odd.mem_bank[1768],db_even.mem_bank[1768]);
$fdisplay(file, "0xDD20,0x%h_0x%h", db_odd.mem_bank[1769],db_even.mem_bank[1769]);
$fdisplay(file, "0xDD40,0x%h_0x%h", db_odd.mem_bank[1770],db_even.mem_bank[1770]);
$fdisplay(file, "0xDD60,0x%h_0x%h", db_odd.mem_bank[1771],db_even.mem_bank[1771]);
$fdisplay(file, "0xDD80,0x%h_0x%h", db_odd.mem_bank[1772],db_even.mem_bank[1772]);
$fdisplay(file, "0xDDA0,0x%h_0x%h", db_odd.mem_bank[1773],db_even.mem_bank[1773]);
$fdisplay(file, "0xDDC0,0x%h_0x%h", db_odd.mem_bank[1774],db_even.mem_bank[1774]);
$fdisplay(file, "0xDDE0,0x%h_0x%h", db_odd.mem_bank[1775],db_even.mem_bank[1775]);
$fdisplay(file, "0xDE00,0x%h_0x%h", db_odd.mem_bank[1776],db_even.mem_bank[1776]);
$fdisplay(file, "0xDE20,0x%h_0x%h", db_odd.mem_bank[1777],db_even.mem_bank[1777]);
$fdisplay(file, "0xDE40,0x%h_0x%h", db_odd.mem_bank[1778],db_even.mem_bank[1778]);
$fdisplay(file, "0xDE60,0x%h_0x%h", db_odd.mem_bank[1779],db_even.mem_bank[1779]);
$fdisplay(file, "0xDE80,0x%h_0x%h", db_odd.mem_bank[1780],db_even.mem_bank[1780]);
$fdisplay(file, "0xDEA0,0x%h_0x%h", db_odd.mem_bank[1781],db_even.mem_bank[1781]);
$fdisplay(file, "0xDEC0,0x%h_0x%h", db_odd.mem_bank[1782],db_even.mem_bank[1782]);
$fdisplay(file, "0xDEE0,0x%h_0x%h", db_odd.mem_bank[1783],db_even.mem_bank[1783]);
$fdisplay(file, "0xDF00,0x%h_0x%h", db_odd.mem_bank[1784],db_even.mem_bank[1784]);
$fdisplay(file, "0xDF20,0x%h_0x%h", db_odd.mem_bank[1785],db_even.mem_bank[1785]);
$fdisplay(file, "0xDF40,0x%h_0x%h", db_odd.mem_bank[1786],db_even.mem_bank[1786]);
$fdisplay(file, "0xDF60,0x%h_0x%h", db_odd.mem_bank[1787],db_even.mem_bank[1787]);
$fdisplay(file, "0xDF80,0x%h_0x%h", db_odd.mem_bank[1788],db_even.mem_bank[1788]);
$fdisplay(file, "0xDFA0,0x%h_0x%h", db_odd.mem_bank[1789],db_even.mem_bank[1789]);
$fdisplay(file, "0xDFC0,0x%h_0x%h", db_odd.mem_bank[1790],db_even.mem_bank[1790]);
$fdisplay(file, "0xDFE0,0x%h_0x%h", db_odd.mem_bank[1791],db_even.mem_bank[1791]);
$fdisplay(file, "0xE000,0x%h_0x%h", db_odd.mem_bank[1792],db_even.mem_bank[1792]);
$fdisplay(file, "0xE020,0x%h_0x%h", db_odd.mem_bank[1793],db_even.mem_bank[1793]);
$fdisplay(file, "0xE040,0x%h_0x%h", db_odd.mem_bank[1794],db_even.mem_bank[1794]);
$fdisplay(file, "0xE060,0x%h_0x%h", db_odd.mem_bank[1795],db_even.mem_bank[1795]);
$fdisplay(file, "0xE080,0x%h_0x%h", db_odd.mem_bank[1796],db_even.mem_bank[1796]);
$fdisplay(file, "0xE0A0,0x%h_0x%h", db_odd.mem_bank[1797],db_even.mem_bank[1797]);
$fdisplay(file, "0xE0C0,0x%h_0x%h", db_odd.mem_bank[1798],db_even.mem_bank[1798]);
$fdisplay(file, "0xE0E0,0x%h_0x%h", db_odd.mem_bank[1799],db_even.mem_bank[1799]);
$fdisplay(file, "0xE100,0x%h_0x%h", db_odd.mem_bank[1800],db_even.mem_bank[1800]);
$fdisplay(file, "0xE120,0x%h_0x%h", db_odd.mem_bank[1801],db_even.mem_bank[1801]);
$fdisplay(file, "0xE140,0x%h_0x%h", db_odd.mem_bank[1802],db_even.mem_bank[1802]);
$fdisplay(file, "0xE160,0x%h_0x%h", db_odd.mem_bank[1803],db_even.mem_bank[1803]);
$fdisplay(file, "0xE180,0x%h_0x%h", db_odd.mem_bank[1804],db_even.mem_bank[1804]);
$fdisplay(file, "0xE1A0,0x%h_0x%h", db_odd.mem_bank[1805],db_even.mem_bank[1805]);
$fdisplay(file, "0xE1C0,0x%h_0x%h", db_odd.mem_bank[1806],db_even.mem_bank[1806]);
$fdisplay(file, "0xE1E0,0x%h_0x%h", db_odd.mem_bank[1807],db_even.mem_bank[1807]);
$fdisplay(file, "0xE200,0x%h_0x%h", db_odd.mem_bank[1808],db_even.mem_bank[1808]);
$fdisplay(file, "0xE220,0x%h_0x%h", db_odd.mem_bank[1809],db_even.mem_bank[1809]);
$fdisplay(file, "0xE240,0x%h_0x%h", db_odd.mem_bank[1810],db_even.mem_bank[1810]);
$fdisplay(file, "0xE260,0x%h_0x%h", db_odd.mem_bank[1811],db_even.mem_bank[1811]);
$fdisplay(file, "0xE280,0x%h_0x%h", db_odd.mem_bank[1812],db_even.mem_bank[1812]);
$fdisplay(file, "0xE2A0,0x%h_0x%h", db_odd.mem_bank[1813],db_even.mem_bank[1813]);
$fdisplay(file, "0xE2C0,0x%h_0x%h", db_odd.mem_bank[1814],db_even.mem_bank[1814]);
$fdisplay(file, "0xE2E0,0x%h_0x%h", db_odd.mem_bank[1815],db_even.mem_bank[1815]);
$fdisplay(file, "0xE300,0x%h_0x%h", db_odd.mem_bank[1816],db_even.mem_bank[1816]);
$fdisplay(file, "0xE320,0x%h_0x%h", db_odd.mem_bank[1817],db_even.mem_bank[1817]);
$fdisplay(file, "0xE340,0x%h_0x%h", db_odd.mem_bank[1818],db_even.mem_bank[1818]);
$fdisplay(file, "0xE360,0x%h_0x%h", db_odd.mem_bank[1819],db_even.mem_bank[1819]);
$fdisplay(file, "0xE380,0x%h_0x%h", db_odd.mem_bank[1820],db_even.mem_bank[1820]);
$fdisplay(file, "0xE3A0,0x%h_0x%h", db_odd.mem_bank[1821],db_even.mem_bank[1821]);
$fdisplay(file, "0xE3C0,0x%h_0x%h", db_odd.mem_bank[1822],db_even.mem_bank[1822]);
$fdisplay(file, "0xE3E0,0x%h_0x%h", db_odd.mem_bank[1823],db_even.mem_bank[1823]);
$fdisplay(file, "0xE400,0x%h_0x%h", db_odd.mem_bank[1824],db_even.mem_bank[1824]);
$fdisplay(file, "0xE420,0x%h_0x%h", db_odd.mem_bank[1825],db_even.mem_bank[1825]);
$fdisplay(file, "0xE440,0x%h_0x%h", db_odd.mem_bank[1826],db_even.mem_bank[1826]);
$fdisplay(file, "0xE460,0x%h_0x%h", db_odd.mem_bank[1827],db_even.mem_bank[1827]);
$fdisplay(file, "0xE480,0x%h_0x%h", db_odd.mem_bank[1828],db_even.mem_bank[1828]);
$fdisplay(file, "0xE4A0,0x%h_0x%h", db_odd.mem_bank[1829],db_even.mem_bank[1829]);
$fdisplay(file, "0xE4C0,0x%h_0x%h", db_odd.mem_bank[1830],db_even.mem_bank[1830]);
$fdisplay(file, "0xE4E0,0x%h_0x%h", db_odd.mem_bank[1831],db_even.mem_bank[1831]);
$fdisplay(file, "0xE500,0x%h_0x%h", db_odd.mem_bank[1832],db_even.mem_bank[1832]);
$fdisplay(file, "0xE520,0x%h_0x%h", db_odd.mem_bank[1833],db_even.mem_bank[1833]);
$fdisplay(file, "0xE540,0x%h_0x%h", db_odd.mem_bank[1834],db_even.mem_bank[1834]);
$fdisplay(file, "0xE560,0x%h_0x%h", db_odd.mem_bank[1835],db_even.mem_bank[1835]);
$fdisplay(file, "0xE580,0x%h_0x%h", db_odd.mem_bank[1836],db_even.mem_bank[1836]);
$fdisplay(file, "0xE5A0,0x%h_0x%h", db_odd.mem_bank[1837],db_even.mem_bank[1837]);
$fdisplay(file, "0xE5C0,0x%h_0x%h", db_odd.mem_bank[1838],db_even.mem_bank[1838]);
$fdisplay(file, "0xE5E0,0x%h_0x%h", db_odd.mem_bank[1839],db_even.mem_bank[1839]);
$fdisplay(file, "0xE600,0x%h_0x%h", db_odd.mem_bank[1840],db_even.mem_bank[1840]);
$fdisplay(file, "0xE620,0x%h_0x%h", db_odd.mem_bank[1841],db_even.mem_bank[1841]);
$fdisplay(file, "0xE640,0x%h_0x%h", db_odd.mem_bank[1842],db_even.mem_bank[1842]);
$fdisplay(file, "0xE660,0x%h_0x%h", db_odd.mem_bank[1843],db_even.mem_bank[1843]);
$fdisplay(file, "0xE680,0x%h_0x%h", db_odd.mem_bank[1844],db_even.mem_bank[1844]);
$fdisplay(file, "0xE6A0,0x%h_0x%h", db_odd.mem_bank[1845],db_even.mem_bank[1845]);
$fdisplay(file, "0xE6C0,0x%h_0x%h", db_odd.mem_bank[1846],db_even.mem_bank[1846]);
$fdisplay(file, "0xE6E0,0x%h_0x%h", db_odd.mem_bank[1847],db_even.mem_bank[1847]);
$fdisplay(file, "0xE700,0x%h_0x%h", db_odd.mem_bank[1848],db_even.mem_bank[1848]);
$fdisplay(file, "0xE720,0x%h_0x%h", db_odd.mem_bank[1849],db_even.mem_bank[1849]);
$fdisplay(file, "0xE740,0x%h_0x%h", db_odd.mem_bank[1850],db_even.mem_bank[1850]);
$fdisplay(file, "0xE760,0x%h_0x%h", db_odd.mem_bank[1851],db_even.mem_bank[1851]);
$fdisplay(file, "0xE780,0x%h_0x%h", db_odd.mem_bank[1852],db_even.mem_bank[1852]);
$fdisplay(file, "0xE7A0,0x%h_0x%h", db_odd.mem_bank[1853],db_even.mem_bank[1853]);
$fdisplay(file, "0xE7C0,0x%h_0x%h", db_odd.mem_bank[1854],db_even.mem_bank[1854]);
$fdisplay(file, "0xE7E0,0x%h_0x%h", db_odd.mem_bank[1855],db_even.mem_bank[1855]);
$fdisplay(file, "0xE800,0x%h_0x%h", db_odd.mem_bank[1856],db_even.mem_bank[1856]);
$fdisplay(file, "0xE820,0x%h_0x%h", db_odd.mem_bank[1857],db_even.mem_bank[1857]);
$fdisplay(file, "0xE840,0x%h_0x%h", db_odd.mem_bank[1858],db_even.mem_bank[1858]);
$fdisplay(file, "0xE860,0x%h_0x%h", db_odd.mem_bank[1859],db_even.mem_bank[1859]);
$fdisplay(file, "0xE880,0x%h_0x%h", db_odd.mem_bank[1860],db_even.mem_bank[1860]);
$fdisplay(file, "0xE8A0,0x%h_0x%h", db_odd.mem_bank[1861],db_even.mem_bank[1861]);
$fdisplay(file, "0xE8C0,0x%h_0x%h", db_odd.mem_bank[1862],db_even.mem_bank[1862]);
$fdisplay(file, "0xE8E0,0x%h_0x%h", db_odd.mem_bank[1863],db_even.mem_bank[1863]);
$fdisplay(file, "0xE900,0x%h_0x%h", db_odd.mem_bank[1864],db_even.mem_bank[1864]);
$fdisplay(file, "0xE920,0x%h_0x%h", db_odd.mem_bank[1865],db_even.mem_bank[1865]);
$fdisplay(file, "0xE940,0x%h_0x%h", db_odd.mem_bank[1866],db_even.mem_bank[1866]);
$fdisplay(file, "0xE960,0x%h_0x%h", db_odd.mem_bank[1867],db_even.mem_bank[1867]);
$fdisplay(file, "0xE980,0x%h_0x%h", db_odd.mem_bank[1868],db_even.mem_bank[1868]);
$fdisplay(file, "0xE9A0,0x%h_0x%h", db_odd.mem_bank[1869],db_even.mem_bank[1869]);
$fdisplay(file, "0xE9C0,0x%h_0x%h", db_odd.mem_bank[1870],db_even.mem_bank[1870]);
$fdisplay(file, "0xE9E0,0x%h_0x%h", db_odd.mem_bank[1871],db_even.mem_bank[1871]);
$fdisplay(file, "0xEA00,0x%h_0x%h", db_odd.mem_bank[1872],db_even.mem_bank[1872]);
$fdisplay(file, "0xEA20,0x%h_0x%h", db_odd.mem_bank[1873],db_even.mem_bank[1873]);
$fdisplay(file, "0xEA40,0x%h_0x%h", db_odd.mem_bank[1874],db_even.mem_bank[1874]);
$fdisplay(file, "0xEA60,0x%h_0x%h", db_odd.mem_bank[1875],db_even.mem_bank[1875]);
$fdisplay(file, "0xEA80,0x%h_0x%h", db_odd.mem_bank[1876],db_even.mem_bank[1876]);
$fdisplay(file, "0xEAA0,0x%h_0x%h", db_odd.mem_bank[1877],db_even.mem_bank[1877]);
$fdisplay(file, "0xEAC0,0x%h_0x%h", db_odd.mem_bank[1878],db_even.mem_bank[1878]);
$fdisplay(file, "0xEAE0,0x%h_0x%h", db_odd.mem_bank[1879],db_even.mem_bank[1879]);
$fdisplay(file, "0xEB00,0x%h_0x%h", db_odd.mem_bank[1880],db_even.mem_bank[1880]);
$fdisplay(file, "0xEB20,0x%h_0x%h", db_odd.mem_bank[1881],db_even.mem_bank[1881]);
$fdisplay(file, "0xEB40,0x%h_0x%h", db_odd.mem_bank[1882],db_even.mem_bank[1882]);
$fdisplay(file, "0xEB60,0x%h_0x%h", db_odd.mem_bank[1883],db_even.mem_bank[1883]);
$fdisplay(file, "0xEB80,0x%h_0x%h", db_odd.mem_bank[1884],db_even.mem_bank[1884]);
$fdisplay(file, "0xEBA0,0x%h_0x%h", db_odd.mem_bank[1885],db_even.mem_bank[1885]);
$fdisplay(file, "0xEBC0,0x%h_0x%h", db_odd.mem_bank[1886],db_even.mem_bank[1886]);
$fdisplay(file, "0xEBE0,0x%h_0x%h", db_odd.mem_bank[1887],db_even.mem_bank[1887]);
$fdisplay(file, "0xEC00,0x%h_0x%h", db_odd.mem_bank[1888],db_even.mem_bank[1888]);
$fdisplay(file, "0xEC20,0x%h_0x%h", db_odd.mem_bank[1889],db_even.mem_bank[1889]);
$fdisplay(file, "0xEC40,0x%h_0x%h", db_odd.mem_bank[1890],db_even.mem_bank[1890]);
$fdisplay(file, "0xEC60,0x%h_0x%h", db_odd.mem_bank[1891],db_even.mem_bank[1891]);
$fdisplay(file, "0xEC80,0x%h_0x%h", db_odd.mem_bank[1892],db_even.mem_bank[1892]);
$fdisplay(file, "0xECA0,0x%h_0x%h", db_odd.mem_bank[1893],db_even.mem_bank[1893]);
$fdisplay(file, "0xECC0,0x%h_0x%h", db_odd.mem_bank[1894],db_even.mem_bank[1894]);
$fdisplay(file, "0xECE0,0x%h_0x%h", db_odd.mem_bank[1895],db_even.mem_bank[1895]);
$fdisplay(file, "0xED00,0x%h_0x%h", db_odd.mem_bank[1896],db_even.mem_bank[1896]);
$fdisplay(file, "0xED20,0x%h_0x%h", db_odd.mem_bank[1897],db_even.mem_bank[1897]);
$fdisplay(file, "0xED40,0x%h_0x%h", db_odd.mem_bank[1898],db_even.mem_bank[1898]);
$fdisplay(file, "0xED60,0x%h_0x%h", db_odd.mem_bank[1899],db_even.mem_bank[1899]);
$fdisplay(file, "0xED80,0x%h_0x%h", db_odd.mem_bank[1900],db_even.mem_bank[1900]);
$fdisplay(file, "0xEDA0,0x%h_0x%h", db_odd.mem_bank[1901],db_even.mem_bank[1901]);
$fdisplay(file, "0xEDC0,0x%h_0x%h", db_odd.mem_bank[1902],db_even.mem_bank[1902]);
$fdisplay(file, "0xEDE0,0x%h_0x%h", db_odd.mem_bank[1903],db_even.mem_bank[1903]);
$fdisplay(file, "0xEE00,0x%h_0x%h", db_odd.mem_bank[1904],db_even.mem_bank[1904]);
$fdisplay(file, "0xEE20,0x%h_0x%h", db_odd.mem_bank[1905],db_even.mem_bank[1905]);
$fdisplay(file, "0xEE40,0x%h_0x%h", db_odd.mem_bank[1906],db_even.mem_bank[1906]);
$fdisplay(file, "0xEE60,0x%h_0x%h", db_odd.mem_bank[1907],db_even.mem_bank[1907]);
$fdisplay(file, "0xEE80,0x%h_0x%h", db_odd.mem_bank[1908],db_even.mem_bank[1908]);
$fdisplay(file, "0xEEA0,0x%h_0x%h", db_odd.mem_bank[1909],db_even.mem_bank[1909]);
$fdisplay(file, "0xEEC0,0x%h_0x%h", db_odd.mem_bank[1910],db_even.mem_bank[1910]);
$fdisplay(file, "0xEEE0,0x%h_0x%h", db_odd.mem_bank[1911],db_even.mem_bank[1911]);
$fdisplay(file, "0xEF00,0x%h_0x%h", db_odd.mem_bank[1912],db_even.mem_bank[1912]);
$fdisplay(file, "0xEF20,0x%h_0x%h", db_odd.mem_bank[1913],db_even.mem_bank[1913]);
$fdisplay(file, "0xEF40,0x%h_0x%h", db_odd.mem_bank[1914],db_even.mem_bank[1914]);
$fdisplay(file, "0xEF60,0x%h_0x%h", db_odd.mem_bank[1915],db_even.mem_bank[1915]);
$fdisplay(file, "0xEF80,0x%h_0x%h", db_odd.mem_bank[1916],db_even.mem_bank[1916]);
$fdisplay(file, "0xEFA0,0x%h_0x%h", db_odd.mem_bank[1917],db_even.mem_bank[1917]);
$fdisplay(file, "0xEFC0,0x%h_0x%h", db_odd.mem_bank[1918],db_even.mem_bank[1918]);
$fdisplay(file, "0xEFE0,0x%h_0x%h", db_odd.mem_bank[1919],db_even.mem_bank[1919]);
$fdisplay(file, "0xF000,0x%h_0x%h", db_odd.mem_bank[1920],db_even.mem_bank[1920]);
$fdisplay(file, "0xF020,0x%h_0x%h", db_odd.mem_bank[1921],db_even.mem_bank[1921]);
$fdisplay(file, "0xF040,0x%h_0x%h", db_odd.mem_bank[1922],db_even.mem_bank[1922]);
$fdisplay(file, "0xF060,0x%h_0x%h", db_odd.mem_bank[1923],db_even.mem_bank[1923]);
$fdisplay(file, "0xF080,0x%h_0x%h", db_odd.mem_bank[1924],db_even.mem_bank[1924]);
$fdisplay(file, "0xF0A0,0x%h_0x%h", db_odd.mem_bank[1925],db_even.mem_bank[1925]);
$fdisplay(file, "0xF0C0,0x%h_0x%h", db_odd.mem_bank[1926],db_even.mem_bank[1926]);
$fdisplay(file, "0xF0E0,0x%h_0x%h", db_odd.mem_bank[1927],db_even.mem_bank[1927]);
$fdisplay(file, "0xF100,0x%h_0x%h", db_odd.mem_bank[1928],db_even.mem_bank[1928]);
$fdisplay(file, "0xF120,0x%h_0x%h", db_odd.mem_bank[1929],db_even.mem_bank[1929]);
$fdisplay(file, "0xF140,0x%h_0x%h", db_odd.mem_bank[1930],db_even.mem_bank[1930]);
$fdisplay(file, "0xF160,0x%h_0x%h", db_odd.mem_bank[1931],db_even.mem_bank[1931]);
$fdisplay(file, "0xF180,0x%h_0x%h", db_odd.mem_bank[1932],db_even.mem_bank[1932]);
$fdisplay(file, "0xF1A0,0x%h_0x%h", db_odd.mem_bank[1933],db_even.mem_bank[1933]);
$fdisplay(file, "0xF1C0,0x%h_0x%h", db_odd.mem_bank[1934],db_even.mem_bank[1934]);
$fdisplay(file, "0xF1E0,0x%h_0x%h", db_odd.mem_bank[1935],db_even.mem_bank[1935]);
$fdisplay(file, "0xF200,0x%h_0x%h", db_odd.mem_bank[1936],db_even.mem_bank[1936]);
$fdisplay(file, "0xF220,0x%h_0x%h", db_odd.mem_bank[1937],db_even.mem_bank[1937]);
$fdisplay(file, "0xF240,0x%h_0x%h", db_odd.mem_bank[1938],db_even.mem_bank[1938]);
$fdisplay(file, "0xF260,0x%h_0x%h", db_odd.mem_bank[1939],db_even.mem_bank[1939]);
$fdisplay(file, "0xF280,0x%h_0x%h", db_odd.mem_bank[1940],db_even.mem_bank[1940]);
$fdisplay(file, "0xF2A0,0x%h_0x%h", db_odd.mem_bank[1941],db_even.mem_bank[1941]);
$fdisplay(file, "0xF2C0,0x%h_0x%h", db_odd.mem_bank[1942],db_even.mem_bank[1942]);
$fdisplay(file, "0xF2E0,0x%h_0x%h", db_odd.mem_bank[1943],db_even.mem_bank[1943]);
$fdisplay(file, "0xF300,0x%h_0x%h", db_odd.mem_bank[1944],db_even.mem_bank[1944]);
$fdisplay(file, "0xF320,0x%h_0x%h", db_odd.mem_bank[1945],db_even.mem_bank[1945]);
$fdisplay(file, "0xF340,0x%h_0x%h", db_odd.mem_bank[1946],db_even.mem_bank[1946]);
$fdisplay(file, "0xF360,0x%h_0x%h", db_odd.mem_bank[1947],db_even.mem_bank[1947]);
$fdisplay(file, "0xF380,0x%h_0x%h", db_odd.mem_bank[1948],db_even.mem_bank[1948]);
$fdisplay(file, "0xF3A0,0x%h_0x%h", db_odd.mem_bank[1949],db_even.mem_bank[1949]);
$fdisplay(file, "0xF3C0,0x%h_0x%h", db_odd.mem_bank[1950],db_even.mem_bank[1950]);
$fdisplay(file, "0xF3E0,0x%h_0x%h", db_odd.mem_bank[1951],db_even.mem_bank[1951]);
$fdisplay(file, "0xF400,0x%h_0x%h", db_odd.mem_bank[1952],db_even.mem_bank[1952]);
$fdisplay(file, "0xF420,0x%h_0x%h", db_odd.mem_bank[1953],db_even.mem_bank[1953]);
$fdisplay(file, "0xF440,0x%h_0x%h", db_odd.mem_bank[1954],db_even.mem_bank[1954]);
$fdisplay(file, "0xF460,0x%h_0x%h", db_odd.mem_bank[1955],db_even.mem_bank[1955]);
$fdisplay(file, "0xF480,0x%h_0x%h", db_odd.mem_bank[1956],db_even.mem_bank[1956]);
$fdisplay(file, "0xF4A0,0x%h_0x%h", db_odd.mem_bank[1957],db_even.mem_bank[1957]);
$fdisplay(file, "0xF4C0,0x%h_0x%h", db_odd.mem_bank[1958],db_even.mem_bank[1958]);
$fdisplay(file, "0xF4E0,0x%h_0x%h", db_odd.mem_bank[1959],db_even.mem_bank[1959]);
$fdisplay(file, "0xF500,0x%h_0x%h", db_odd.mem_bank[1960],db_even.mem_bank[1960]);
$fdisplay(file, "0xF520,0x%h_0x%h", db_odd.mem_bank[1961],db_even.mem_bank[1961]);
$fdisplay(file, "0xF540,0x%h_0x%h", db_odd.mem_bank[1962],db_even.mem_bank[1962]);
$fdisplay(file, "0xF560,0x%h_0x%h", db_odd.mem_bank[1963],db_even.mem_bank[1963]);
$fdisplay(file, "0xF580,0x%h_0x%h", db_odd.mem_bank[1964],db_even.mem_bank[1964]);
$fdisplay(file, "0xF5A0,0x%h_0x%h", db_odd.mem_bank[1965],db_even.mem_bank[1965]);
$fdisplay(file, "0xF5C0,0x%h_0x%h", db_odd.mem_bank[1966],db_even.mem_bank[1966]);
$fdisplay(file, "0xF5E0,0x%h_0x%h", db_odd.mem_bank[1967],db_even.mem_bank[1967]);
$fdisplay(file, "0xF600,0x%h_0x%h", db_odd.mem_bank[1968],db_even.mem_bank[1968]);
$fdisplay(file, "0xF620,0x%h_0x%h", db_odd.mem_bank[1969],db_even.mem_bank[1969]);
$fdisplay(file, "0xF640,0x%h_0x%h", db_odd.mem_bank[1970],db_even.mem_bank[1970]);
$fdisplay(file, "0xF660,0x%h_0x%h", db_odd.mem_bank[1971],db_even.mem_bank[1971]);
$fdisplay(file, "0xF680,0x%h_0x%h", db_odd.mem_bank[1972],db_even.mem_bank[1972]);
$fdisplay(file, "0xF6A0,0x%h_0x%h", db_odd.mem_bank[1973],db_even.mem_bank[1973]);
$fdisplay(file, "0xF6C0,0x%h_0x%h", db_odd.mem_bank[1974],db_even.mem_bank[1974]);
$fdisplay(file, "0xF6E0,0x%h_0x%h", db_odd.mem_bank[1975],db_even.mem_bank[1975]);
$fdisplay(file, "0xF700,0x%h_0x%h", db_odd.mem_bank[1976],db_even.mem_bank[1976]);
$fdisplay(file, "0xF720,0x%h_0x%h", db_odd.mem_bank[1977],db_even.mem_bank[1977]);
$fdisplay(file, "0xF740,0x%h_0x%h", db_odd.mem_bank[1978],db_even.mem_bank[1978]);
$fdisplay(file, "0xF760,0x%h_0x%h", db_odd.mem_bank[1979],db_even.mem_bank[1979]);
$fdisplay(file, "0xF780,0x%h_0x%h", db_odd.mem_bank[1980],db_even.mem_bank[1980]);
$fdisplay(file, "0xF7A0,0x%h_0x%h", db_odd.mem_bank[1981],db_even.mem_bank[1981]);
$fdisplay(file, "0xF7C0,0x%h_0x%h", db_odd.mem_bank[1982],db_even.mem_bank[1982]);
$fdisplay(file, "0xF7E0,0x%h_0x%h", db_odd.mem_bank[1983],db_even.mem_bank[1983]);
$fdisplay(file, "0xF800,0x%h_0x%h", db_odd.mem_bank[1984],db_even.mem_bank[1984]);
$fdisplay(file, "0xF820,0x%h_0x%h", db_odd.mem_bank[1985],db_even.mem_bank[1985]);
$fdisplay(file, "0xF840,0x%h_0x%h", db_odd.mem_bank[1986],db_even.mem_bank[1986]);
$fdisplay(file, "0xF860,0x%h_0x%h", db_odd.mem_bank[1987],db_even.mem_bank[1987]);
$fdisplay(file, "0xF880,0x%h_0x%h", db_odd.mem_bank[1988],db_even.mem_bank[1988]);
$fdisplay(file, "0xF8A0,0x%h_0x%h", db_odd.mem_bank[1989],db_even.mem_bank[1989]);
$fdisplay(file, "0xF8C0,0x%h_0x%h", db_odd.mem_bank[1990],db_even.mem_bank[1990]);
$fdisplay(file, "0xF8E0,0x%h_0x%h", db_odd.mem_bank[1991],db_even.mem_bank[1991]);
$fdisplay(file, "0xF900,0x%h_0x%h", db_odd.mem_bank[1992],db_even.mem_bank[1992]);
$fdisplay(file, "0xF920,0x%h_0x%h", db_odd.mem_bank[1993],db_even.mem_bank[1993]);
$fdisplay(file, "0xF940,0x%h_0x%h", db_odd.mem_bank[1994],db_even.mem_bank[1994]);
$fdisplay(file, "0xF960,0x%h_0x%h", db_odd.mem_bank[1995],db_even.mem_bank[1995]);
$fdisplay(file, "0xF980,0x%h_0x%h", db_odd.mem_bank[1996],db_even.mem_bank[1996]);
$fdisplay(file, "0xF9A0,0x%h_0x%h", db_odd.mem_bank[1997],db_even.mem_bank[1997]);
$fdisplay(file, "0xF9C0,0x%h_0x%h", db_odd.mem_bank[1998],db_even.mem_bank[1998]);
$fdisplay(file, "0xF9E0,0x%h_0x%h", db_odd.mem_bank[1999],db_even.mem_bank[1999]);
$fdisplay(file, "0xFA00,0x%h_0x%h", db_odd.mem_bank[2000],db_even.mem_bank[2000]);
$fdisplay(file, "0xFA20,0x%h_0x%h", db_odd.mem_bank[2001],db_even.mem_bank[2001]);
$fdisplay(file, "0xFA40,0x%h_0x%h", db_odd.mem_bank[2002],db_even.mem_bank[2002]);
$fdisplay(file, "0xFA60,0x%h_0x%h", db_odd.mem_bank[2003],db_even.mem_bank[2003]);
$fdisplay(file, "0xFA80,0x%h_0x%h", db_odd.mem_bank[2004],db_even.mem_bank[2004]);
$fdisplay(file, "0xFAA0,0x%h_0x%h", db_odd.mem_bank[2005],db_even.mem_bank[2005]);
$fdisplay(file, "0xFAC0,0x%h_0x%h", db_odd.mem_bank[2006],db_even.mem_bank[2006]);
$fdisplay(file, "0xFAE0,0x%h_0x%h", db_odd.mem_bank[2007],db_even.mem_bank[2007]);
$fdisplay(file, "0xFB00,0x%h_0x%h", db_odd.mem_bank[2008],db_even.mem_bank[2008]);
$fdisplay(file, "0xFB20,0x%h_0x%h", db_odd.mem_bank[2009],db_even.mem_bank[2009]);
$fdisplay(file, "0xFB40,0x%h_0x%h", db_odd.mem_bank[2010],db_even.mem_bank[2010]);
$fdisplay(file, "0xFB60,0x%h_0x%h", db_odd.mem_bank[2011],db_even.mem_bank[2011]);
$fdisplay(file, "0xFB80,0x%h_0x%h", db_odd.mem_bank[2012],db_even.mem_bank[2012]);
$fdisplay(file, "0xFBA0,0x%h_0x%h", db_odd.mem_bank[2013],db_even.mem_bank[2013]);
$fdisplay(file, "0xFBC0,0x%h_0x%h", db_odd.mem_bank[2014],db_even.mem_bank[2014]);
$fdisplay(file, "0xFBE0,0x%h_0x%h", db_odd.mem_bank[2015],db_even.mem_bank[2015]);
$fdisplay(file, "0xFC00,0x%h_0x%h", db_odd.mem_bank[2016],db_even.mem_bank[2016]);
$fdisplay(file, "0xFC20,0x%h_0x%h", db_odd.mem_bank[2017],db_even.mem_bank[2017]);
$fdisplay(file, "0xFC40,0x%h_0x%h", db_odd.mem_bank[2018],db_even.mem_bank[2018]);
$fdisplay(file, "0xFC60,0x%h_0x%h", db_odd.mem_bank[2019],db_even.mem_bank[2019]);
$fdisplay(file, "0xFC80,0x%h_0x%h", db_odd.mem_bank[2020],db_even.mem_bank[2020]);
$fdisplay(file, "0xFCA0,0x%h_0x%h", db_odd.mem_bank[2021],db_even.mem_bank[2021]);
$fdisplay(file, "0xFCC0,0x%h_0x%h", db_odd.mem_bank[2022],db_even.mem_bank[2022]);
$fdisplay(file, "0xFCE0,0x%h_0x%h", db_odd.mem_bank[2023],db_even.mem_bank[2023]);
$fdisplay(file, "0xFD00,0x%h_0x%h", db_odd.mem_bank[2024],db_even.mem_bank[2024]);
$fdisplay(file, "0xFD20,0x%h_0x%h", db_odd.mem_bank[2025],db_even.mem_bank[2025]);
$fdisplay(file, "0xFD40,0x%h_0x%h", db_odd.mem_bank[2026],db_even.mem_bank[2026]);
$fdisplay(file, "0xFD60,0x%h_0x%h", db_odd.mem_bank[2027],db_even.mem_bank[2027]);
$fdisplay(file, "0xFD80,0x%h_0x%h", db_odd.mem_bank[2028],db_even.mem_bank[2028]);
$fdisplay(file, "0xFDA0,0x%h_0x%h", db_odd.mem_bank[2029],db_even.mem_bank[2029]);
$fdisplay(file, "0xFDC0,0x%h_0x%h", db_odd.mem_bank[2030],db_even.mem_bank[2030]);
$fdisplay(file, "0xFDE0,0x%h_0x%h", db_odd.mem_bank[2031],db_even.mem_bank[2031]);
$fdisplay(file, "0xFE00,0x%h_0x%h", db_odd.mem_bank[2032],db_even.mem_bank[2032]);
$fdisplay(file, "0xFE20,0x%h_0x%h", db_odd.mem_bank[2033],db_even.mem_bank[2033]);
$fdisplay(file, "0xFE40,0x%h_0x%h", db_odd.mem_bank[2034],db_even.mem_bank[2034]);
$fdisplay(file, "0xFE60,0x%h_0x%h", db_odd.mem_bank[2035],db_even.mem_bank[2035]);
$fdisplay(file, "0xFE80,0x%h_0x%h", db_odd.mem_bank[2036],db_even.mem_bank[2036]);
$fdisplay(file, "0xFEA0,0x%h_0x%h", db_odd.mem_bank[2037],db_even.mem_bank[2037]);
$fdisplay(file, "0xFEC0,0x%h_0x%h", db_odd.mem_bank[2038],db_even.mem_bank[2038]);
$fdisplay(file, "0xFEE0,0x%h_0x%h", db_odd.mem_bank[2039],db_even.mem_bank[2039]);
$fdisplay(file, "0xFF00,0x%h_0x%h", db_odd.mem_bank[2040],db_even.mem_bank[2040]);
$fdisplay(file, "0xFF20,0x%h_0x%h", db_odd.mem_bank[2041],db_even.mem_bank[2041]);
$fdisplay(file, "0xFF40,0x%h_0x%h", db_odd.mem_bank[2042],db_even.mem_bank[2042]);
$fdisplay(file, "0xFF60,0x%h_0x%h", db_odd.mem_bank[2043],db_even.mem_bank[2043]);
$fdisplay(file, "0xFF80,0x%h_0x%h", db_odd.mem_bank[2044],db_even.mem_bank[2044]);
$fdisplay(file, "0xFFA0,0x%h_0x%h", db_odd.mem_bank[2045],db_even.mem_bank[2045]);
$fdisplay(file, "0xFFC0,0x%h_0x%h", db_odd.mem_bank[2046],db_even.mem_bank[2046]);
$fdisplay(file, "0xFFE0,0x%h_0x%h", db_odd.mem_bank[2047],db_even.mem_bank[2047]);
$fdisplay(file, "0x10000,0x%h_0x%h", db_odd.mem_bank[2048],db_even.mem_bank[2048]);
$fdisplay(file, "0x10020,0x%h_0x%h", db_odd.mem_bank[2049],db_even.mem_bank[2049]);
$fdisplay(file, "0x10040,0x%h_0x%h", db_odd.mem_bank[2050],db_even.mem_bank[2050]);
$fdisplay(file, "0x10060,0x%h_0x%h", db_odd.mem_bank[2051],db_even.mem_bank[2051]);
$fdisplay(file, "0x10080,0x%h_0x%h", db_odd.mem_bank[2052],db_even.mem_bank[2052]);
$fdisplay(file, "0x100A0,0x%h_0x%h", db_odd.mem_bank[2053],db_even.mem_bank[2053]);
$fdisplay(file, "0x100C0,0x%h_0x%h", db_odd.mem_bank[2054],db_even.mem_bank[2054]);
$fdisplay(file, "0x100E0,0x%h_0x%h", db_odd.mem_bank[2055],db_even.mem_bank[2055]);
$fdisplay(file, "0x10100,0x%h_0x%h", db_odd.mem_bank[2056],db_even.mem_bank[2056]);
$fdisplay(file, "0x10120,0x%h_0x%h", db_odd.mem_bank[2057],db_even.mem_bank[2057]);
$fdisplay(file, "0x10140,0x%h_0x%h", db_odd.mem_bank[2058],db_even.mem_bank[2058]);
$fdisplay(file, "0x10160,0x%h_0x%h", db_odd.mem_bank[2059],db_even.mem_bank[2059]);
$fdisplay(file, "0x10180,0x%h_0x%h", db_odd.mem_bank[2060],db_even.mem_bank[2060]);
$fdisplay(file, "0x101A0,0x%h_0x%h", db_odd.mem_bank[2061],db_even.mem_bank[2061]);
$fdisplay(file, "0x101C0,0x%h_0x%h", db_odd.mem_bank[2062],db_even.mem_bank[2062]);
$fdisplay(file, "0x101E0,0x%h_0x%h", db_odd.mem_bank[2063],db_even.mem_bank[2063]);
$fdisplay(file, "0x10200,0x%h_0x%h", db_odd.mem_bank[2064],db_even.mem_bank[2064]);
$fdisplay(file, "0x10220,0x%h_0x%h", db_odd.mem_bank[2065],db_even.mem_bank[2065]);
$fdisplay(file, "0x10240,0x%h_0x%h", db_odd.mem_bank[2066],db_even.mem_bank[2066]);
$fdisplay(file, "0x10260,0x%h_0x%h", db_odd.mem_bank[2067],db_even.mem_bank[2067]);
$fdisplay(file, "0x10280,0x%h_0x%h", db_odd.mem_bank[2068],db_even.mem_bank[2068]);
$fdisplay(file, "0x102A0,0x%h_0x%h", db_odd.mem_bank[2069],db_even.mem_bank[2069]);
$fdisplay(file, "0x102C0,0x%h_0x%h", db_odd.mem_bank[2070],db_even.mem_bank[2070]);
$fdisplay(file, "0x102E0,0x%h_0x%h", db_odd.mem_bank[2071],db_even.mem_bank[2071]);
$fdisplay(file, "0x10300,0x%h_0x%h", db_odd.mem_bank[2072],db_even.mem_bank[2072]);
$fdisplay(file, "0x10320,0x%h_0x%h", db_odd.mem_bank[2073],db_even.mem_bank[2073]);
$fdisplay(file, "0x10340,0x%h_0x%h", db_odd.mem_bank[2074],db_even.mem_bank[2074]);
$fdisplay(file, "0x10360,0x%h_0x%h", db_odd.mem_bank[2075],db_even.mem_bank[2075]);
$fdisplay(file, "0x10380,0x%h_0x%h", db_odd.mem_bank[2076],db_even.mem_bank[2076]);
$fdisplay(file, "0x103A0,0x%h_0x%h", db_odd.mem_bank[2077],db_even.mem_bank[2077]);
$fdisplay(file, "0x103C0,0x%h_0x%h", db_odd.mem_bank[2078],db_even.mem_bank[2078]);
$fdisplay(file, "0x103E0,0x%h_0x%h", db_odd.mem_bank[2079],db_even.mem_bank[2079]);
$fdisplay(file, "0x10400,0x%h_0x%h", db_odd.mem_bank[2080],db_even.mem_bank[2080]);
$fdisplay(file, "0x10420,0x%h_0x%h", db_odd.mem_bank[2081],db_even.mem_bank[2081]);
$fdisplay(file, "0x10440,0x%h_0x%h", db_odd.mem_bank[2082],db_even.mem_bank[2082]);
$fdisplay(file, "0x10460,0x%h_0x%h", db_odd.mem_bank[2083],db_even.mem_bank[2083]);
$fdisplay(file, "0x10480,0x%h_0x%h", db_odd.mem_bank[2084],db_even.mem_bank[2084]);
$fdisplay(file, "0x104A0,0x%h_0x%h", db_odd.mem_bank[2085],db_even.mem_bank[2085]);
$fdisplay(file, "0x104C0,0x%h_0x%h", db_odd.mem_bank[2086],db_even.mem_bank[2086]);
$fdisplay(file, "0x104E0,0x%h_0x%h", db_odd.mem_bank[2087],db_even.mem_bank[2087]);
$fdisplay(file, "0x10500,0x%h_0x%h", db_odd.mem_bank[2088],db_even.mem_bank[2088]);
$fdisplay(file, "0x10520,0x%h_0x%h", db_odd.mem_bank[2089],db_even.mem_bank[2089]);
$fdisplay(file, "0x10540,0x%h_0x%h", db_odd.mem_bank[2090],db_even.mem_bank[2090]);
$fdisplay(file, "0x10560,0x%h_0x%h", db_odd.mem_bank[2091],db_even.mem_bank[2091]);
$fdisplay(file, "0x10580,0x%h_0x%h", db_odd.mem_bank[2092],db_even.mem_bank[2092]);
$fdisplay(file, "0x105A0,0x%h_0x%h", db_odd.mem_bank[2093],db_even.mem_bank[2093]);
$fdisplay(file, "0x105C0,0x%h_0x%h", db_odd.mem_bank[2094],db_even.mem_bank[2094]);
$fdisplay(file, "0x105E0,0x%h_0x%h", db_odd.mem_bank[2095],db_even.mem_bank[2095]);
$fdisplay(file, "0x10600,0x%h_0x%h", db_odd.mem_bank[2096],db_even.mem_bank[2096]);
$fdisplay(file, "0x10620,0x%h_0x%h", db_odd.mem_bank[2097],db_even.mem_bank[2097]);
$fdisplay(file, "0x10640,0x%h_0x%h", db_odd.mem_bank[2098],db_even.mem_bank[2098]);
$fdisplay(file, "0x10660,0x%h_0x%h", db_odd.mem_bank[2099],db_even.mem_bank[2099]);
$fdisplay(file, "0x10680,0x%h_0x%h", db_odd.mem_bank[2100],db_even.mem_bank[2100]);
$fdisplay(file, "0x106A0,0x%h_0x%h", db_odd.mem_bank[2101],db_even.mem_bank[2101]);
$fdisplay(file, "0x106C0,0x%h_0x%h", db_odd.mem_bank[2102],db_even.mem_bank[2102]);
$fdisplay(file, "0x106E0,0x%h_0x%h", db_odd.mem_bank[2103],db_even.mem_bank[2103]);
$fdisplay(file, "0x10700,0x%h_0x%h", db_odd.mem_bank[2104],db_even.mem_bank[2104]);
$fdisplay(file, "0x10720,0x%h_0x%h", db_odd.mem_bank[2105],db_even.mem_bank[2105]);
$fdisplay(file, "0x10740,0x%h_0x%h", db_odd.mem_bank[2106],db_even.mem_bank[2106]);
$fdisplay(file, "0x10760,0x%h_0x%h", db_odd.mem_bank[2107],db_even.mem_bank[2107]);
$fdisplay(file, "0x10780,0x%h_0x%h", db_odd.mem_bank[2108],db_even.mem_bank[2108]);
$fdisplay(file, "0x107A0,0x%h_0x%h", db_odd.mem_bank[2109],db_even.mem_bank[2109]);
$fdisplay(file, "0x107C0,0x%h_0x%h", db_odd.mem_bank[2110],db_even.mem_bank[2110]);
$fdisplay(file, "0x107E0,0x%h_0x%h", db_odd.mem_bank[2111],db_even.mem_bank[2111]);
$fdisplay(file, "0x10800,0x%h_0x%h", db_odd.mem_bank[2112],db_even.mem_bank[2112]);
$fdisplay(file, "0x10820,0x%h_0x%h", db_odd.mem_bank[2113],db_even.mem_bank[2113]);
$fdisplay(file, "0x10840,0x%h_0x%h", db_odd.mem_bank[2114],db_even.mem_bank[2114]);
$fdisplay(file, "0x10860,0x%h_0x%h", db_odd.mem_bank[2115],db_even.mem_bank[2115]);
$fdisplay(file, "0x10880,0x%h_0x%h", db_odd.mem_bank[2116],db_even.mem_bank[2116]);
$fdisplay(file, "0x108A0,0x%h_0x%h", db_odd.mem_bank[2117],db_even.mem_bank[2117]);
$fdisplay(file, "0x108C0,0x%h_0x%h", db_odd.mem_bank[2118],db_even.mem_bank[2118]);
$fdisplay(file, "0x108E0,0x%h_0x%h", db_odd.mem_bank[2119],db_even.mem_bank[2119]);
$fdisplay(file, "0x10900,0x%h_0x%h", db_odd.mem_bank[2120],db_even.mem_bank[2120]);
$fdisplay(file, "0x10920,0x%h_0x%h", db_odd.mem_bank[2121],db_even.mem_bank[2121]);
$fdisplay(file, "0x10940,0x%h_0x%h", db_odd.mem_bank[2122],db_even.mem_bank[2122]);
$fdisplay(file, "0x10960,0x%h_0x%h", db_odd.mem_bank[2123],db_even.mem_bank[2123]);
$fdisplay(file, "0x10980,0x%h_0x%h", db_odd.mem_bank[2124],db_even.mem_bank[2124]);
$fdisplay(file, "0x109A0,0x%h_0x%h", db_odd.mem_bank[2125],db_even.mem_bank[2125]);
$fdisplay(file, "0x109C0,0x%h_0x%h", db_odd.mem_bank[2126],db_even.mem_bank[2126]);
$fdisplay(file, "0x109E0,0x%h_0x%h", db_odd.mem_bank[2127],db_even.mem_bank[2127]);
$fdisplay(file, "0x10A00,0x%h_0x%h", db_odd.mem_bank[2128],db_even.mem_bank[2128]);
$fdisplay(file, "0x10A20,0x%h_0x%h", db_odd.mem_bank[2129],db_even.mem_bank[2129]);
$fdisplay(file, "0x10A40,0x%h_0x%h", db_odd.mem_bank[2130],db_even.mem_bank[2130]);
$fdisplay(file, "0x10A60,0x%h_0x%h", db_odd.mem_bank[2131],db_even.mem_bank[2131]);
$fdisplay(file, "0x10A80,0x%h_0x%h", db_odd.mem_bank[2132],db_even.mem_bank[2132]);
$fdisplay(file, "0x10AA0,0x%h_0x%h", db_odd.mem_bank[2133],db_even.mem_bank[2133]);
$fdisplay(file, "0x10AC0,0x%h_0x%h", db_odd.mem_bank[2134],db_even.mem_bank[2134]);
$fdisplay(file, "0x10AE0,0x%h_0x%h", db_odd.mem_bank[2135],db_even.mem_bank[2135]);
$fdisplay(file, "0x10B00,0x%h_0x%h", db_odd.mem_bank[2136],db_even.mem_bank[2136]);
$fdisplay(file, "0x10B20,0x%h_0x%h", db_odd.mem_bank[2137],db_even.mem_bank[2137]);
$fdisplay(file, "0x10B40,0x%h_0x%h", db_odd.mem_bank[2138],db_even.mem_bank[2138]);
$fdisplay(file, "0x10B60,0x%h_0x%h", db_odd.mem_bank[2139],db_even.mem_bank[2139]);
$fdisplay(file, "0x10B80,0x%h_0x%h", db_odd.mem_bank[2140],db_even.mem_bank[2140]);
$fdisplay(file, "0x10BA0,0x%h_0x%h", db_odd.mem_bank[2141],db_even.mem_bank[2141]);
$fdisplay(file, "0x10BC0,0x%h_0x%h", db_odd.mem_bank[2142],db_even.mem_bank[2142]);
$fdisplay(file, "0x10BE0,0x%h_0x%h", db_odd.mem_bank[2143],db_even.mem_bank[2143]);
$fdisplay(file, "0x10C00,0x%h_0x%h", db_odd.mem_bank[2144],db_even.mem_bank[2144]);
$fdisplay(file, "0x10C20,0x%h_0x%h", db_odd.mem_bank[2145],db_even.mem_bank[2145]);
$fdisplay(file, "0x10C40,0x%h_0x%h", db_odd.mem_bank[2146],db_even.mem_bank[2146]);
$fdisplay(file, "0x10C60,0x%h_0x%h", db_odd.mem_bank[2147],db_even.mem_bank[2147]);
$fdisplay(file, "0x10C80,0x%h_0x%h", db_odd.mem_bank[2148],db_even.mem_bank[2148]);
$fdisplay(file, "0x10CA0,0x%h_0x%h", db_odd.mem_bank[2149],db_even.mem_bank[2149]);
$fdisplay(file, "0x10CC0,0x%h_0x%h", db_odd.mem_bank[2150],db_even.mem_bank[2150]);
$fdisplay(file, "0x10CE0,0x%h_0x%h", db_odd.mem_bank[2151],db_even.mem_bank[2151]);
$fdisplay(file, "0x10D00,0x%h_0x%h", db_odd.mem_bank[2152],db_even.mem_bank[2152]);
$fdisplay(file, "0x10D20,0x%h_0x%h", db_odd.mem_bank[2153],db_even.mem_bank[2153]);
$fdisplay(file, "0x10D40,0x%h_0x%h", db_odd.mem_bank[2154],db_even.mem_bank[2154]);
$fdisplay(file, "0x10D60,0x%h_0x%h", db_odd.mem_bank[2155],db_even.mem_bank[2155]);
$fdisplay(file, "0x10D80,0x%h_0x%h", db_odd.mem_bank[2156],db_even.mem_bank[2156]);
$fdisplay(file, "0x10DA0,0x%h_0x%h", db_odd.mem_bank[2157],db_even.mem_bank[2157]);
$fdisplay(file, "0x10DC0,0x%h_0x%h", db_odd.mem_bank[2158],db_even.mem_bank[2158]);
$fdisplay(file, "0x10DE0,0x%h_0x%h", db_odd.mem_bank[2159],db_even.mem_bank[2159]);
$fdisplay(file, "0x10E00,0x%h_0x%h", db_odd.mem_bank[2160],db_even.mem_bank[2160]);
$fdisplay(file, "0x10E20,0x%h_0x%h", db_odd.mem_bank[2161],db_even.mem_bank[2161]);
$fdisplay(file, "0x10E40,0x%h_0x%h", db_odd.mem_bank[2162],db_even.mem_bank[2162]);
$fdisplay(file, "0x10E60,0x%h_0x%h", db_odd.mem_bank[2163],db_even.mem_bank[2163]);
$fdisplay(file, "0x10E80,0x%h_0x%h", db_odd.mem_bank[2164],db_even.mem_bank[2164]);
$fdisplay(file, "0x10EA0,0x%h_0x%h", db_odd.mem_bank[2165],db_even.mem_bank[2165]);
$fdisplay(file, "0x10EC0,0x%h_0x%h", db_odd.mem_bank[2166],db_even.mem_bank[2166]);
$fdisplay(file, "0x10EE0,0x%h_0x%h", db_odd.mem_bank[2167],db_even.mem_bank[2167]);
$fdisplay(file, "0x10F00,0x%h_0x%h", db_odd.mem_bank[2168],db_even.mem_bank[2168]);
$fdisplay(file, "0x10F20,0x%h_0x%h", db_odd.mem_bank[2169],db_even.mem_bank[2169]);
$fdisplay(file, "0x10F40,0x%h_0x%h", db_odd.mem_bank[2170],db_even.mem_bank[2170]);
$fdisplay(file, "0x10F60,0x%h_0x%h", db_odd.mem_bank[2171],db_even.mem_bank[2171]);
$fdisplay(file, "0x10F80,0x%h_0x%h", db_odd.mem_bank[2172],db_even.mem_bank[2172]);
$fdisplay(file, "0x10FA0,0x%h_0x%h", db_odd.mem_bank[2173],db_even.mem_bank[2173]);
$fdisplay(file, "0x10FC0,0x%h_0x%h", db_odd.mem_bank[2174],db_even.mem_bank[2174]);
$fdisplay(file, "0x10FE0,0x%h_0x%h", db_odd.mem_bank[2175],db_even.mem_bank[2175]);
$fdisplay(file, "0x11000,0x%h_0x%h", db_odd.mem_bank[2176],db_even.mem_bank[2176]);
$fdisplay(file, "0x11020,0x%h_0x%h", db_odd.mem_bank[2177],db_even.mem_bank[2177]);
$fdisplay(file, "0x11040,0x%h_0x%h", db_odd.mem_bank[2178],db_even.mem_bank[2178]);
$fdisplay(file, "0x11060,0x%h_0x%h", db_odd.mem_bank[2179],db_even.mem_bank[2179]);
$fdisplay(file, "0x11080,0x%h_0x%h", db_odd.mem_bank[2180],db_even.mem_bank[2180]);
$fdisplay(file, "0x110A0,0x%h_0x%h", db_odd.mem_bank[2181],db_even.mem_bank[2181]);
$fdisplay(file, "0x110C0,0x%h_0x%h", db_odd.mem_bank[2182],db_even.mem_bank[2182]);
$fdisplay(file, "0x110E0,0x%h_0x%h", db_odd.mem_bank[2183],db_even.mem_bank[2183]);
$fdisplay(file, "0x11100,0x%h_0x%h", db_odd.mem_bank[2184],db_even.mem_bank[2184]);
$fdisplay(file, "0x11120,0x%h_0x%h", db_odd.mem_bank[2185],db_even.mem_bank[2185]);
$fdisplay(file, "0x11140,0x%h_0x%h", db_odd.mem_bank[2186],db_even.mem_bank[2186]);
$fdisplay(file, "0x11160,0x%h_0x%h", db_odd.mem_bank[2187],db_even.mem_bank[2187]);
$fdisplay(file, "0x11180,0x%h_0x%h", db_odd.mem_bank[2188],db_even.mem_bank[2188]);
$fdisplay(file, "0x111A0,0x%h_0x%h", db_odd.mem_bank[2189],db_even.mem_bank[2189]);
$fdisplay(file, "0x111C0,0x%h_0x%h", db_odd.mem_bank[2190],db_even.mem_bank[2190]);
$fdisplay(file, "0x111E0,0x%h_0x%h", db_odd.mem_bank[2191],db_even.mem_bank[2191]);
$fdisplay(file, "0x11200,0x%h_0x%h", db_odd.mem_bank[2192],db_even.mem_bank[2192]);
$fdisplay(file, "0x11220,0x%h_0x%h", db_odd.mem_bank[2193],db_even.mem_bank[2193]);
$fdisplay(file, "0x11240,0x%h_0x%h", db_odd.mem_bank[2194],db_even.mem_bank[2194]);
$fdisplay(file, "0x11260,0x%h_0x%h", db_odd.mem_bank[2195],db_even.mem_bank[2195]);
$fdisplay(file, "0x11280,0x%h_0x%h", db_odd.mem_bank[2196],db_even.mem_bank[2196]);
$fdisplay(file, "0x112A0,0x%h_0x%h", db_odd.mem_bank[2197],db_even.mem_bank[2197]);
$fdisplay(file, "0x112C0,0x%h_0x%h", db_odd.mem_bank[2198],db_even.mem_bank[2198]);
$fdisplay(file, "0x112E0,0x%h_0x%h", db_odd.mem_bank[2199],db_even.mem_bank[2199]);
$fdisplay(file, "0x11300,0x%h_0x%h", db_odd.mem_bank[2200],db_even.mem_bank[2200]);
$fdisplay(file, "0x11320,0x%h_0x%h", db_odd.mem_bank[2201],db_even.mem_bank[2201]);
$fdisplay(file, "0x11340,0x%h_0x%h", db_odd.mem_bank[2202],db_even.mem_bank[2202]);
$fdisplay(file, "0x11360,0x%h_0x%h", db_odd.mem_bank[2203],db_even.mem_bank[2203]);
$fdisplay(file, "0x11380,0x%h_0x%h", db_odd.mem_bank[2204],db_even.mem_bank[2204]);
$fdisplay(file, "0x113A0,0x%h_0x%h", db_odd.mem_bank[2205],db_even.mem_bank[2205]);
$fdisplay(file, "0x113C0,0x%h_0x%h", db_odd.mem_bank[2206],db_even.mem_bank[2206]);
$fdisplay(file, "0x113E0,0x%h_0x%h", db_odd.mem_bank[2207],db_even.mem_bank[2207]);
$fdisplay(file, "0x11400,0x%h_0x%h", db_odd.mem_bank[2208],db_even.mem_bank[2208]);
$fdisplay(file, "0x11420,0x%h_0x%h", db_odd.mem_bank[2209],db_even.mem_bank[2209]);
$fdisplay(file, "0x11440,0x%h_0x%h", db_odd.mem_bank[2210],db_even.mem_bank[2210]);
$fdisplay(file, "0x11460,0x%h_0x%h", db_odd.mem_bank[2211],db_even.mem_bank[2211]);
$fdisplay(file, "0x11480,0x%h_0x%h", db_odd.mem_bank[2212],db_even.mem_bank[2212]);
$fdisplay(file, "0x114A0,0x%h_0x%h", db_odd.mem_bank[2213],db_even.mem_bank[2213]);
$fdisplay(file, "0x114C0,0x%h_0x%h", db_odd.mem_bank[2214],db_even.mem_bank[2214]);
$fdisplay(file, "0x114E0,0x%h_0x%h", db_odd.mem_bank[2215],db_even.mem_bank[2215]);
$fdisplay(file, "0x11500,0x%h_0x%h", db_odd.mem_bank[2216],db_even.mem_bank[2216]);
$fdisplay(file, "0x11520,0x%h_0x%h", db_odd.mem_bank[2217],db_even.mem_bank[2217]);
$fdisplay(file, "0x11540,0x%h_0x%h", db_odd.mem_bank[2218],db_even.mem_bank[2218]);
$fdisplay(file, "0x11560,0x%h_0x%h", db_odd.mem_bank[2219],db_even.mem_bank[2219]);
$fdisplay(file, "0x11580,0x%h_0x%h", db_odd.mem_bank[2220],db_even.mem_bank[2220]);
$fdisplay(file, "0x115A0,0x%h_0x%h", db_odd.mem_bank[2221],db_even.mem_bank[2221]);
$fdisplay(file, "0x115C0,0x%h_0x%h", db_odd.mem_bank[2222],db_even.mem_bank[2222]);
$fdisplay(file, "0x115E0,0x%h_0x%h", db_odd.mem_bank[2223],db_even.mem_bank[2223]);
$fdisplay(file, "0x11600,0x%h_0x%h", db_odd.mem_bank[2224],db_even.mem_bank[2224]);
$fdisplay(file, "0x11620,0x%h_0x%h", db_odd.mem_bank[2225],db_even.mem_bank[2225]);
$fdisplay(file, "0x11640,0x%h_0x%h", db_odd.mem_bank[2226],db_even.mem_bank[2226]);
$fdisplay(file, "0x11660,0x%h_0x%h", db_odd.mem_bank[2227],db_even.mem_bank[2227]);
$fdisplay(file, "0x11680,0x%h_0x%h", db_odd.mem_bank[2228],db_even.mem_bank[2228]);
$fdisplay(file, "0x116A0,0x%h_0x%h", db_odd.mem_bank[2229],db_even.mem_bank[2229]);
$fdisplay(file, "0x116C0,0x%h_0x%h", db_odd.mem_bank[2230],db_even.mem_bank[2230]);
$fdisplay(file, "0x116E0,0x%h_0x%h", db_odd.mem_bank[2231],db_even.mem_bank[2231]);
$fdisplay(file, "0x11700,0x%h_0x%h", db_odd.mem_bank[2232],db_even.mem_bank[2232]);
$fdisplay(file, "0x11720,0x%h_0x%h", db_odd.mem_bank[2233],db_even.mem_bank[2233]);
$fdisplay(file, "0x11740,0x%h_0x%h", db_odd.mem_bank[2234],db_even.mem_bank[2234]);
$fdisplay(file, "0x11760,0x%h_0x%h", db_odd.mem_bank[2235],db_even.mem_bank[2235]);
$fdisplay(file, "0x11780,0x%h_0x%h", db_odd.mem_bank[2236],db_even.mem_bank[2236]);
$fdisplay(file, "0x117A0,0x%h_0x%h", db_odd.mem_bank[2237],db_even.mem_bank[2237]);
$fdisplay(file, "0x117C0,0x%h_0x%h", db_odd.mem_bank[2238],db_even.mem_bank[2238]);
$fdisplay(file, "0x117E0,0x%h_0x%h", db_odd.mem_bank[2239],db_even.mem_bank[2239]);
$fdisplay(file, "0x11800,0x%h_0x%h", db_odd.mem_bank[2240],db_even.mem_bank[2240]);
$fdisplay(file, "0x11820,0x%h_0x%h", db_odd.mem_bank[2241],db_even.mem_bank[2241]);
$fdisplay(file, "0x11840,0x%h_0x%h", db_odd.mem_bank[2242],db_even.mem_bank[2242]);
$fdisplay(file, "0x11860,0x%h_0x%h", db_odd.mem_bank[2243],db_even.mem_bank[2243]);
$fdisplay(file, "0x11880,0x%h_0x%h", db_odd.mem_bank[2244],db_even.mem_bank[2244]);
$fdisplay(file, "0x118A0,0x%h_0x%h", db_odd.mem_bank[2245],db_even.mem_bank[2245]);
$fdisplay(file, "0x118C0,0x%h_0x%h", db_odd.mem_bank[2246],db_even.mem_bank[2246]);
$fdisplay(file, "0x118E0,0x%h_0x%h", db_odd.mem_bank[2247],db_even.mem_bank[2247]);
$fdisplay(file, "0x11900,0x%h_0x%h", db_odd.mem_bank[2248],db_even.mem_bank[2248]);
$fdisplay(file, "0x11920,0x%h_0x%h", db_odd.mem_bank[2249],db_even.mem_bank[2249]);
$fdisplay(file, "0x11940,0x%h_0x%h", db_odd.mem_bank[2250],db_even.mem_bank[2250]);
$fdisplay(file, "0x11960,0x%h_0x%h", db_odd.mem_bank[2251],db_even.mem_bank[2251]);
$fdisplay(file, "0x11980,0x%h_0x%h", db_odd.mem_bank[2252],db_even.mem_bank[2252]);
$fdisplay(file, "0x119A0,0x%h_0x%h", db_odd.mem_bank[2253],db_even.mem_bank[2253]);
$fdisplay(file, "0x119C0,0x%h_0x%h", db_odd.mem_bank[2254],db_even.mem_bank[2254]);
$fdisplay(file, "0x119E0,0x%h_0x%h", db_odd.mem_bank[2255],db_even.mem_bank[2255]);
$fdisplay(file, "0x11A00,0x%h_0x%h", db_odd.mem_bank[2256],db_even.mem_bank[2256]);
$fdisplay(file, "0x11A20,0x%h_0x%h", db_odd.mem_bank[2257],db_even.mem_bank[2257]);
$fdisplay(file, "0x11A40,0x%h_0x%h", db_odd.mem_bank[2258],db_even.mem_bank[2258]);
$fdisplay(file, "0x11A60,0x%h_0x%h", db_odd.mem_bank[2259],db_even.mem_bank[2259]);
$fdisplay(file, "0x11A80,0x%h_0x%h", db_odd.mem_bank[2260],db_even.mem_bank[2260]);
$fdisplay(file, "0x11AA0,0x%h_0x%h", db_odd.mem_bank[2261],db_even.mem_bank[2261]);
$fdisplay(file, "0x11AC0,0x%h_0x%h", db_odd.mem_bank[2262],db_even.mem_bank[2262]);
$fdisplay(file, "0x11AE0,0x%h_0x%h", db_odd.mem_bank[2263],db_even.mem_bank[2263]);
$fdisplay(file, "0x11B00,0x%h_0x%h", db_odd.mem_bank[2264],db_even.mem_bank[2264]);
$fdisplay(file, "0x11B20,0x%h_0x%h", db_odd.mem_bank[2265],db_even.mem_bank[2265]);
$fdisplay(file, "0x11B40,0x%h_0x%h", db_odd.mem_bank[2266],db_even.mem_bank[2266]);
$fdisplay(file, "0x11B60,0x%h_0x%h", db_odd.mem_bank[2267],db_even.mem_bank[2267]);
$fdisplay(file, "0x11B80,0x%h_0x%h", db_odd.mem_bank[2268],db_even.mem_bank[2268]);
$fdisplay(file, "0x11BA0,0x%h_0x%h", db_odd.mem_bank[2269],db_even.mem_bank[2269]);
$fdisplay(file, "0x11BC0,0x%h_0x%h", db_odd.mem_bank[2270],db_even.mem_bank[2270]);
$fdisplay(file, "0x11BE0,0x%h_0x%h", db_odd.mem_bank[2271],db_even.mem_bank[2271]);
$fdisplay(file, "0x11C00,0x%h_0x%h", db_odd.mem_bank[2272],db_even.mem_bank[2272]);
$fdisplay(file, "0x11C20,0x%h_0x%h", db_odd.mem_bank[2273],db_even.mem_bank[2273]);
$fdisplay(file, "0x11C40,0x%h_0x%h", db_odd.mem_bank[2274],db_even.mem_bank[2274]);
$fdisplay(file, "0x11C60,0x%h_0x%h", db_odd.mem_bank[2275],db_even.mem_bank[2275]);
$fdisplay(file, "0x11C80,0x%h_0x%h", db_odd.mem_bank[2276],db_even.mem_bank[2276]);
$fdisplay(file, "0x11CA0,0x%h_0x%h", db_odd.mem_bank[2277],db_even.mem_bank[2277]);
$fdisplay(file, "0x11CC0,0x%h_0x%h", db_odd.mem_bank[2278],db_even.mem_bank[2278]);
$fdisplay(file, "0x11CE0,0x%h_0x%h", db_odd.mem_bank[2279],db_even.mem_bank[2279]);
$fdisplay(file, "0x11D00,0x%h_0x%h", db_odd.mem_bank[2280],db_even.mem_bank[2280]);
$fdisplay(file, "0x11D20,0x%h_0x%h", db_odd.mem_bank[2281],db_even.mem_bank[2281]);
$fdisplay(file, "0x11D40,0x%h_0x%h", db_odd.mem_bank[2282],db_even.mem_bank[2282]);
$fdisplay(file, "0x11D60,0x%h_0x%h", db_odd.mem_bank[2283],db_even.mem_bank[2283]);
$fdisplay(file, "0x11D80,0x%h_0x%h", db_odd.mem_bank[2284],db_even.mem_bank[2284]);
$fdisplay(file, "0x11DA0,0x%h_0x%h", db_odd.mem_bank[2285],db_even.mem_bank[2285]);
$fdisplay(file, "0x11DC0,0x%h_0x%h", db_odd.mem_bank[2286],db_even.mem_bank[2286]);
$fdisplay(file, "0x11DE0,0x%h_0x%h", db_odd.mem_bank[2287],db_even.mem_bank[2287]);
$fdisplay(file, "0x11E00,0x%h_0x%h", db_odd.mem_bank[2288],db_even.mem_bank[2288]);
$fdisplay(file, "0x11E20,0x%h_0x%h", db_odd.mem_bank[2289],db_even.mem_bank[2289]);
$fdisplay(file, "0x11E40,0x%h_0x%h", db_odd.mem_bank[2290],db_even.mem_bank[2290]);
$fdisplay(file, "0x11E60,0x%h_0x%h", db_odd.mem_bank[2291],db_even.mem_bank[2291]);
$fdisplay(file, "0x11E80,0x%h_0x%h", db_odd.mem_bank[2292],db_even.mem_bank[2292]);
$fdisplay(file, "0x11EA0,0x%h_0x%h", db_odd.mem_bank[2293],db_even.mem_bank[2293]);
$fdisplay(file, "0x11EC0,0x%h_0x%h", db_odd.mem_bank[2294],db_even.mem_bank[2294]);
$fdisplay(file, "0x11EE0,0x%h_0x%h", db_odd.mem_bank[2295],db_even.mem_bank[2295]);
$fdisplay(file, "0x11F00,0x%h_0x%h", db_odd.mem_bank[2296],db_even.mem_bank[2296]);
$fdisplay(file, "0x11F20,0x%h_0x%h", db_odd.mem_bank[2297],db_even.mem_bank[2297]);
$fdisplay(file, "0x11F40,0x%h_0x%h", db_odd.mem_bank[2298],db_even.mem_bank[2298]);
$fdisplay(file, "0x11F60,0x%h_0x%h", db_odd.mem_bank[2299],db_even.mem_bank[2299]);
$fdisplay(file, "0x11F80,0x%h_0x%h", db_odd.mem_bank[2300],db_even.mem_bank[2300]);
$fdisplay(file, "0x11FA0,0x%h_0x%h", db_odd.mem_bank[2301],db_even.mem_bank[2301]);
$fdisplay(file, "0x11FC0,0x%h_0x%h", db_odd.mem_bank[2302],db_even.mem_bank[2302]);
$fdisplay(file, "0x11FE0,0x%h_0x%h", db_odd.mem_bank[2303],db_even.mem_bank[2303]);
$fdisplay(file, "0x12000,0x%h_0x%h", db_odd.mem_bank[2304],db_even.mem_bank[2304]);
$fdisplay(file, "0x12020,0x%h_0x%h", db_odd.mem_bank[2305],db_even.mem_bank[2305]);
$fdisplay(file, "0x12040,0x%h_0x%h", db_odd.mem_bank[2306],db_even.mem_bank[2306]);
$fdisplay(file, "0x12060,0x%h_0x%h", db_odd.mem_bank[2307],db_even.mem_bank[2307]);
$fdisplay(file, "0x12080,0x%h_0x%h", db_odd.mem_bank[2308],db_even.mem_bank[2308]);
$fdisplay(file, "0x120A0,0x%h_0x%h", db_odd.mem_bank[2309],db_even.mem_bank[2309]);
$fdisplay(file, "0x120C0,0x%h_0x%h", db_odd.mem_bank[2310],db_even.mem_bank[2310]);
$fdisplay(file, "0x120E0,0x%h_0x%h", db_odd.mem_bank[2311],db_even.mem_bank[2311]);
$fdisplay(file, "0x12100,0x%h_0x%h", db_odd.mem_bank[2312],db_even.mem_bank[2312]);
$fdisplay(file, "0x12120,0x%h_0x%h", db_odd.mem_bank[2313],db_even.mem_bank[2313]);
$fdisplay(file, "0x12140,0x%h_0x%h", db_odd.mem_bank[2314],db_even.mem_bank[2314]);
$fdisplay(file, "0x12160,0x%h_0x%h", db_odd.mem_bank[2315],db_even.mem_bank[2315]);
$fdisplay(file, "0x12180,0x%h_0x%h", db_odd.mem_bank[2316],db_even.mem_bank[2316]);
$fdisplay(file, "0x121A0,0x%h_0x%h", db_odd.mem_bank[2317],db_even.mem_bank[2317]);
$fdisplay(file, "0x121C0,0x%h_0x%h", db_odd.mem_bank[2318],db_even.mem_bank[2318]);
$fdisplay(file, "0x121E0,0x%h_0x%h", db_odd.mem_bank[2319],db_even.mem_bank[2319]);
$fdisplay(file, "0x12200,0x%h_0x%h", db_odd.mem_bank[2320],db_even.mem_bank[2320]);
$fdisplay(file, "0x12220,0x%h_0x%h", db_odd.mem_bank[2321],db_even.mem_bank[2321]);
$fdisplay(file, "0x12240,0x%h_0x%h", db_odd.mem_bank[2322],db_even.mem_bank[2322]);
$fdisplay(file, "0x12260,0x%h_0x%h", db_odd.mem_bank[2323],db_even.mem_bank[2323]);
$fdisplay(file, "0x12280,0x%h_0x%h", db_odd.mem_bank[2324],db_even.mem_bank[2324]);
$fdisplay(file, "0x122A0,0x%h_0x%h", db_odd.mem_bank[2325],db_even.mem_bank[2325]);
$fdisplay(file, "0x122C0,0x%h_0x%h", db_odd.mem_bank[2326],db_even.mem_bank[2326]);
$fdisplay(file, "0x122E0,0x%h_0x%h", db_odd.mem_bank[2327],db_even.mem_bank[2327]);
$fdisplay(file, "0x12300,0x%h_0x%h", db_odd.mem_bank[2328],db_even.mem_bank[2328]);
$fdisplay(file, "0x12320,0x%h_0x%h", db_odd.mem_bank[2329],db_even.mem_bank[2329]);
$fdisplay(file, "0x12340,0x%h_0x%h", db_odd.mem_bank[2330],db_even.mem_bank[2330]);
$fdisplay(file, "0x12360,0x%h_0x%h", db_odd.mem_bank[2331],db_even.mem_bank[2331]);
$fdisplay(file, "0x12380,0x%h_0x%h", db_odd.mem_bank[2332],db_even.mem_bank[2332]);
$fdisplay(file, "0x123A0,0x%h_0x%h", db_odd.mem_bank[2333],db_even.mem_bank[2333]);
$fdisplay(file, "0x123C0,0x%h_0x%h", db_odd.mem_bank[2334],db_even.mem_bank[2334]);
$fdisplay(file, "0x123E0,0x%h_0x%h", db_odd.mem_bank[2335],db_even.mem_bank[2335]);
$fdisplay(file, "0x12400,0x%h_0x%h", db_odd.mem_bank[2336],db_even.mem_bank[2336]);
$fdisplay(file, "0x12420,0x%h_0x%h", db_odd.mem_bank[2337],db_even.mem_bank[2337]);
$fdisplay(file, "0x12440,0x%h_0x%h", db_odd.mem_bank[2338],db_even.mem_bank[2338]);
$fdisplay(file, "0x12460,0x%h_0x%h", db_odd.mem_bank[2339],db_even.mem_bank[2339]);
$fdisplay(file, "0x12480,0x%h_0x%h", db_odd.mem_bank[2340],db_even.mem_bank[2340]);
$fdisplay(file, "0x124A0,0x%h_0x%h", db_odd.mem_bank[2341],db_even.mem_bank[2341]);
$fdisplay(file, "0x124C0,0x%h_0x%h", db_odd.mem_bank[2342],db_even.mem_bank[2342]);
$fdisplay(file, "0x124E0,0x%h_0x%h", db_odd.mem_bank[2343],db_even.mem_bank[2343]);
$fdisplay(file, "0x12500,0x%h_0x%h", db_odd.mem_bank[2344],db_even.mem_bank[2344]);
$fdisplay(file, "0x12520,0x%h_0x%h", db_odd.mem_bank[2345],db_even.mem_bank[2345]);
$fdisplay(file, "0x12540,0x%h_0x%h", db_odd.mem_bank[2346],db_even.mem_bank[2346]);
$fdisplay(file, "0x12560,0x%h_0x%h", db_odd.mem_bank[2347],db_even.mem_bank[2347]);
$fdisplay(file, "0x12580,0x%h_0x%h", db_odd.mem_bank[2348],db_even.mem_bank[2348]);
$fdisplay(file, "0x125A0,0x%h_0x%h", db_odd.mem_bank[2349],db_even.mem_bank[2349]);
$fdisplay(file, "0x125C0,0x%h_0x%h", db_odd.mem_bank[2350],db_even.mem_bank[2350]);
$fdisplay(file, "0x125E0,0x%h_0x%h", db_odd.mem_bank[2351],db_even.mem_bank[2351]);
$fdisplay(file, "0x12600,0x%h_0x%h", db_odd.mem_bank[2352],db_even.mem_bank[2352]);
$fdisplay(file, "0x12620,0x%h_0x%h", db_odd.mem_bank[2353],db_even.mem_bank[2353]);
$fdisplay(file, "0x12640,0x%h_0x%h", db_odd.mem_bank[2354],db_even.mem_bank[2354]);
$fdisplay(file, "0x12660,0x%h_0x%h", db_odd.mem_bank[2355],db_even.mem_bank[2355]);
$fdisplay(file, "0x12680,0x%h_0x%h", db_odd.mem_bank[2356],db_even.mem_bank[2356]);
$fdisplay(file, "0x126A0,0x%h_0x%h", db_odd.mem_bank[2357],db_even.mem_bank[2357]);
$fdisplay(file, "0x126C0,0x%h_0x%h", db_odd.mem_bank[2358],db_even.mem_bank[2358]);
$fdisplay(file, "0x126E0,0x%h_0x%h", db_odd.mem_bank[2359],db_even.mem_bank[2359]);
$fdisplay(file, "0x12700,0x%h_0x%h", db_odd.mem_bank[2360],db_even.mem_bank[2360]);
$fdisplay(file, "0x12720,0x%h_0x%h", db_odd.mem_bank[2361],db_even.mem_bank[2361]);
$fdisplay(file, "0x12740,0x%h_0x%h", db_odd.mem_bank[2362],db_even.mem_bank[2362]);
$fdisplay(file, "0x12760,0x%h_0x%h", db_odd.mem_bank[2363],db_even.mem_bank[2363]);
$fdisplay(file, "0x12780,0x%h_0x%h", db_odd.mem_bank[2364],db_even.mem_bank[2364]);
$fdisplay(file, "0x127A0,0x%h_0x%h", db_odd.mem_bank[2365],db_even.mem_bank[2365]);
$fdisplay(file, "0x127C0,0x%h_0x%h", db_odd.mem_bank[2366],db_even.mem_bank[2366]);
$fdisplay(file, "0x127E0,0x%h_0x%h", db_odd.mem_bank[2367],db_even.mem_bank[2367]);
$fdisplay(file, "0x12800,0x%h_0x%h", db_odd.mem_bank[2368],db_even.mem_bank[2368]);
$fdisplay(file, "0x12820,0x%h_0x%h", db_odd.mem_bank[2369],db_even.mem_bank[2369]);
$fdisplay(file, "0x12840,0x%h_0x%h", db_odd.mem_bank[2370],db_even.mem_bank[2370]);
$fdisplay(file, "0x12860,0x%h_0x%h", db_odd.mem_bank[2371],db_even.mem_bank[2371]);
$fdisplay(file, "0x12880,0x%h_0x%h", db_odd.mem_bank[2372],db_even.mem_bank[2372]);
$fdisplay(file, "0x128A0,0x%h_0x%h", db_odd.mem_bank[2373],db_even.mem_bank[2373]);
$fdisplay(file, "0x128C0,0x%h_0x%h", db_odd.mem_bank[2374],db_even.mem_bank[2374]);
$fdisplay(file, "0x128E0,0x%h_0x%h", db_odd.mem_bank[2375],db_even.mem_bank[2375]);
$fdisplay(file, "0x12900,0x%h_0x%h", db_odd.mem_bank[2376],db_even.mem_bank[2376]);
$fdisplay(file, "0x12920,0x%h_0x%h", db_odd.mem_bank[2377],db_even.mem_bank[2377]);
$fdisplay(file, "0x12940,0x%h_0x%h", db_odd.mem_bank[2378],db_even.mem_bank[2378]);
$fdisplay(file, "0x12960,0x%h_0x%h", db_odd.mem_bank[2379],db_even.mem_bank[2379]);
$fdisplay(file, "0x12980,0x%h_0x%h", db_odd.mem_bank[2380],db_even.mem_bank[2380]);
$fdisplay(file, "0x129A0,0x%h_0x%h", db_odd.mem_bank[2381],db_even.mem_bank[2381]);
$fdisplay(file, "0x129C0,0x%h_0x%h", db_odd.mem_bank[2382],db_even.mem_bank[2382]);
$fdisplay(file, "0x129E0,0x%h_0x%h", db_odd.mem_bank[2383],db_even.mem_bank[2383]);
$fdisplay(file, "0x12A00,0x%h_0x%h", db_odd.mem_bank[2384],db_even.mem_bank[2384]);
$fdisplay(file, "0x12A20,0x%h_0x%h", db_odd.mem_bank[2385],db_even.mem_bank[2385]);
$fdisplay(file, "0x12A40,0x%h_0x%h", db_odd.mem_bank[2386],db_even.mem_bank[2386]);
$fdisplay(file, "0x12A60,0x%h_0x%h", db_odd.mem_bank[2387],db_even.mem_bank[2387]);
$fdisplay(file, "0x12A80,0x%h_0x%h", db_odd.mem_bank[2388],db_even.mem_bank[2388]);
$fdisplay(file, "0x12AA0,0x%h_0x%h", db_odd.mem_bank[2389],db_even.mem_bank[2389]);
$fdisplay(file, "0x12AC0,0x%h_0x%h", db_odd.mem_bank[2390],db_even.mem_bank[2390]);
$fdisplay(file, "0x12AE0,0x%h_0x%h", db_odd.mem_bank[2391],db_even.mem_bank[2391]);
$fdisplay(file, "0x12B00,0x%h_0x%h", db_odd.mem_bank[2392],db_even.mem_bank[2392]);
$fdisplay(file, "0x12B20,0x%h_0x%h", db_odd.mem_bank[2393],db_even.mem_bank[2393]);
$fdisplay(file, "0x12B40,0x%h_0x%h", db_odd.mem_bank[2394],db_even.mem_bank[2394]);
$fdisplay(file, "0x12B60,0x%h_0x%h", db_odd.mem_bank[2395],db_even.mem_bank[2395]);
$fdisplay(file, "0x12B80,0x%h_0x%h", db_odd.mem_bank[2396],db_even.mem_bank[2396]);
$fdisplay(file, "0x12BA0,0x%h_0x%h", db_odd.mem_bank[2397],db_even.mem_bank[2397]);
$fdisplay(file, "0x12BC0,0x%h_0x%h", db_odd.mem_bank[2398],db_even.mem_bank[2398]);
$fdisplay(file, "0x12BE0,0x%h_0x%h", db_odd.mem_bank[2399],db_even.mem_bank[2399]);
$fdisplay(file, "0x12C00,0x%h_0x%h", db_odd.mem_bank[2400],db_even.mem_bank[2400]);
$fdisplay(file, "0x12C20,0x%h_0x%h", db_odd.mem_bank[2401],db_even.mem_bank[2401]);
$fdisplay(file, "0x12C40,0x%h_0x%h", db_odd.mem_bank[2402],db_even.mem_bank[2402]);
$fdisplay(file, "0x12C60,0x%h_0x%h", db_odd.mem_bank[2403],db_even.mem_bank[2403]);
$fdisplay(file, "0x12C80,0x%h_0x%h", db_odd.mem_bank[2404],db_even.mem_bank[2404]);
$fdisplay(file, "0x12CA0,0x%h_0x%h", db_odd.mem_bank[2405],db_even.mem_bank[2405]);
$fdisplay(file, "0x12CC0,0x%h_0x%h", db_odd.mem_bank[2406],db_even.mem_bank[2406]);
$fdisplay(file, "0x12CE0,0x%h_0x%h", db_odd.mem_bank[2407],db_even.mem_bank[2407]);
$fdisplay(file, "0x12D00,0x%h_0x%h", db_odd.mem_bank[2408],db_even.mem_bank[2408]);
$fdisplay(file, "0x12D20,0x%h_0x%h", db_odd.mem_bank[2409],db_even.mem_bank[2409]);
$fdisplay(file, "0x12D40,0x%h_0x%h", db_odd.mem_bank[2410],db_even.mem_bank[2410]);
$fdisplay(file, "0x12D60,0x%h_0x%h", db_odd.mem_bank[2411],db_even.mem_bank[2411]);
$fdisplay(file, "0x12D80,0x%h_0x%h", db_odd.mem_bank[2412],db_even.mem_bank[2412]);
$fdisplay(file, "0x12DA0,0x%h_0x%h", db_odd.mem_bank[2413],db_even.mem_bank[2413]);
$fdisplay(file, "0x12DC0,0x%h_0x%h", db_odd.mem_bank[2414],db_even.mem_bank[2414]);
$fdisplay(file, "0x12DE0,0x%h_0x%h", db_odd.mem_bank[2415],db_even.mem_bank[2415]);
$fdisplay(file, "0x12E00,0x%h_0x%h", db_odd.mem_bank[2416],db_even.mem_bank[2416]);
$fdisplay(file, "0x12E20,0x%h_0x%h", db_odd.mem_bank[2417],db_even.mem_bank[2417]);
$fdisplay(file, "0x12E40,0x%h_0x%h", db_odd.mem_bank[2418],db_even.mem_bank[2418]);
$fdisplay(file, "0x12E60,0x%h_0x%h", db_odd.mem_bank[2419],db_even.mem_bank[2419]);
$fdisplay(file, "0x12E80,0x%h_0x%h", db_odd.mem_bank[2420],db_even.mem_bank[2420]);
$fdisplay(file, "0x12EA0,0x%h_0x%h", db_odd.mem_bank[2421],db_even.mem_bank[2421]);
$fdisplay(file, "0x12EC0,0x%h_0x%h", db_odd.mem_bank[2422],db_even.mem_bank[2422]);
$fdisplay(file, "0x12EE0,0x%h_0x%h", db_odd.mem_bank[2423],db_even.mem_bank[2423]);
$fdisplay(file, "0x12F00,0x%h_0x%h", db_odd.mem_bank[2424],db_even.mem_bank[2424]);
$fdisplay(file, "0x12F20,0x%h_0x%h", db_odd.mem_bank[2425],db_even.mem_bank[2425]);
$fdisplay(file, "0x12F40,0x%h_0x%h", db_odd.mem_bank[2426],db_even.mem_bank[2426]);
$fdisplay(file, "0x12F60,0x%h_0x%h", db_odd.mem_bank[2427],db_even.mem_bank[2427]);
$fdisplay(file, "0x12F80,0x%h_0x%h", db_odd.mem_bank[2428],db_even.mem_bank[2428]);
$fdisplay(file, "0x12FA0,0x%h_0x%h", db_odd.mem_bank[2429],db_even.mem_bank[2429]);
$fdisplay(file, "0x12FC0,0x%h_0x%h", db_odd.mem_bank[2430],db_even.mem_bank[2430]);
$fdisplay(file, "0x12FE0,0x%h_0x%h", db_odd.mem_bank[2431],db_even.mem_bank[2431]);
$fdisplay(file, "0x13000,0x%h_0x%h", db_odd.mem_bank[2432],db_even.mem_bank[2432]);
$fdisplay(file, "0x13020,0x%h_0x%h", db_odd.mem_bank[2433],db_even.mem_bank[2433]);
$fdisplay(file, "0x13040,0x%h_0x%h", db_odd.mem_bank[2434],db_even.mem_bank[2434]);
$fdisplay(file, "0x13060,0x%h_0x%h", db_odd.mem_bank[2435],db_even.mem_bank[2435]);
$fdisplay(file, "0x13080,0x%h_0x%h", db_odd.mem_bank[2436],db_even.mem_bank[2436]);
$fdisplay(file, "0x130A0,0x%h_0x%h", db_odd.mem_bank[2437],db_even.mem_bank[2437]);
$fdisplay(file, "0x130C0,0x%h_0x%h", db_odd.mem_bank[2438],db_even.mem_bank[2438]);
$fdisplay(file, "0x130E0,0x%h_0x%h", db_odd.mem_bank[2439],db_even.mem_bank[2439]);
$fdisplay(file, "0x13100,0x%h_0x%h", db_odd.mem_bank[2440],db_even.mem_bank[2440]);
$fdisplay(file, "0x13120,0x%h_0x%h", db_odd.mem_bank[2441],db_even.mem_bank[2441]);
$fdisplay(file, "0x13140,0x%h_0x%h", db_odd.mem_bank[2442],db_even.mem_bank[2442]);
$fdisplay(file, "0x13160,0x%h_0x%h", db_odd.mem_bank[2443],db_even.mem_bank[2443]);
$fdisplay(file, "0x13180,0x%h_0x%h", db_odd.mem_bank[2444],db_even.mem_bank[2444]);
$fdisplay(file, "0x131A0,0x%h_0x%h", db_odd.mem_bank[2445],db_even.mem_bank[2445]);
$fdisplay(file, "0x131C0,0x%h_0x%h", db_odd.mem_bank[2446],db_even.mem_bank[2446]);
$fdisplay(file, "0x131E0,0x%h_0x%h", db_odd.mem_bank[2447],db_even.mem_bank[2447]);
$fdisplay(file, "0x13200,0x%h_0x%h", db_odd.mem_bank[2448],db_even.mem_bank[2448]);
$fdisplay(file, "0x13220,0x%h_0x%h", db_odd.mem_bank[2449],db_even.mem_bank[2449]);
$fdisplay(file, "0x13240,0x%h_0x%h", db_odd.mem_bank[2450],db_even.mem_bank[2450]);
$fdisplay(file, "0x13260,0x%h_0x%h", db_odd.mem_bank[2451],db_even.mem_bank[2451]);
$fdisplay(file, "0x13280,0x%h_0x%h", db_odd.mem_bank[2452],db_even.mem_bank[2452]);
$fdisplay(file, "0x132A0,0x%h_0x%h", db_odd.mem_bank[2453],db_even.mem_bank[2453]);
$fdisplay(file, "0x132C0,0x%h_0x%h", db_odd.mem_bank[2454],db_even.mem_bank[2454]);
$fdisplay(file, "0x132E0,0x%h_0x%h", db_odd.mem_bank[2455],db_even.mem_bank[2455]);
$fdisplay(file, "0x13300,0x%h_0x%h", db_odd.mem_bank[2456],db_even.mem_bank[2456]);
$fdisplay(file, "0x13320,0x%h_0x%h", db_odd.mem_bank[2457],db_even.mem_bank[2457]);
$fdisplay(file, "0x13340,0x%h_0x%h", db_odd.mem_bank[2458],db_even.mem_bank[2458]);
$fdisplay(file, "0x13360,0x%h_0x%h", db_odd.mem_bank[2459],db_even.mem_bank[2459]);
$fdisplay(file, "0x13380,0x%h_0x%h", db_odd.mem_bank[2460],db_even.mem_bank[2460]);
$fdisplay(file, "0x133A0,0x%h_0x%h", db_odd.mem_bank[2461],db_even.mem_bank[2461]);
$fdisplay(file, "0x133C0,0x%h_0x%h", db_odd.mem_bank[2462],db_even.mem_bank[2462]);
$fdisplay(file, "0x133E0,0x%h_0x%h", db_odd.mem_bank[2463],db_even.mem_bank[2463]);
$fdisplay(file, "0x13400,0x%h_0x%h", db_odd.mem_bank[2464],db_even.mem_bank[2464]);
$fdisplay(file, "0x13420,0x%h_0x%h", db_odd.mem_bank[2465],db_even.mem_bank[2465]);
$fdisplay(file, "0x13440,0x%h_0x%h", db_odd.mem_bank[2466],db_even.mem_bank[2466]);
$fdisplay(file, "0x13460,0x%h_0x%h", db_odd.mem_bank[2467],db_even.mem_bank[2467]);
$fdisplay(file, "0x13480,0x%h_0x%h", db_odd.mem_bank[2468],db_even.mem_bank[2468]);
$fdisplay(file, "0x134A0,0x%h_0x%h", db_odd.mem_bank[2469],db_even.mem_bank[2469]);
$fdisplay(file, "0x134C0,0x%h_0x%h", db_odd.mem_bank[2470],db_even.mem_bank[2470]);
$fdisplay(file, "0x134E0,0x%h_0x%h", db_odd.mem_bank[2471],db_even.mem_bank[2471]);
$fdisplay(file, "0x13500,0x%h_0x%h", db_odd.mem_bank[2472],db_even.mem_bank[2472]);
$fdisplay(file, "0x13520,0x%h_0x%h", db_odd.mem_bank[2473],db_even.mem_bank[2473]);
$fdisplay(file, "0x13540,0x%h_0x%h", db_odd.mem_bank[2474],db_even.mem_bank[2474]);
$fdisplay(file, "0x13560,0x%h_0x%h", db_odd.mem_bank[2475],db_even.mem_bank[2475]);
$fdisplay(file, "0x13580,0x%h_0x%h", db_odd.mem_bank[2476],db_even.mem_bank[2476]);
$fdisplay(file, "0x135A0,0x%h_0x%h", db_odd.mem_bank[2477],db_even.mem_bank[2477]);
$fdisplay(file, "0x135C0,0x%h_0x%h", db_odd.mem_bank[2478],db_even.mem_bank[2478]);
$fdisplay(file, "0x135E0,0x%h_0x%h", db_odd.mem_bank[2479],db_even.mem_bank[2479]);
$fdisplay(file, "0x13600,0x%h_0x%h", db_odd.mem_bank[2480],db_even.mem_bank[2480]);
$fdisplay(file, "0x13620,0x%h_0x%h", db_odd.mem_bank[2481],db_even.mem_bank[2481]);
$fdisplay(file, "0x13640,0x%h_0x%h", db_odd.mem_bank[2482],db_even.mem_bank[2482]);
$fdisplay(file, "0x13660,0x%h_0x%h", db_odd.mem_bank[2483],db_even.mem_bank[2483]);
$fdisplay(file, "0x13680,0x%h_0x%h", db_odd.mem_bank[2484],db_even.mem_bank[2484]);
$fdisplay(file, "0x136A0,0x%h_0x%h", db_odd.mem_bank[2485],db_even.mem_bank[2485]);
$fdisplay(file, "0x136C0,0x%h_0x%h", db_odd.mem_bank[2486],db_even.mem_bank[2486]);
$fdisplay(file, "0x136E0,0x%h_0x%h", db_odd.mem_bank[2487],db_even.mem_bank[2487]);
$fdisplay(file, "0x13700,0x%h_0x%h", db_odd.mem_bank[2488],db_even.mem_bank[2488]);
$fdisplay(file, "0x13720,0x%h_0x%h", db_odd.mem_bank[2489],db_even.mem_bank[2489]);
$fdisplay(file, "0x13740,0x%h_0x%h", db_odd.mem_bank[2490],db_even.mem_bank[2490]);
$fdisplay(file, "0x13760,0x%h_0x%h", db_odd.mem_bank[2491],db_even.mem_bank[2491]);
$fdisplay(file, "0x13780,0x%h_0x%h", db_odd.mem_bank[2492],db_even.mem_bank[2492]);
$fdisplay(file, "0x137A0,0x%h_0x%h", db_odd.mem_bank[2493],db_even.mem_bank[2493]);
$fdisplay(file, "0x137C0,0x%h_0x%h", db_odd.mem_bank[2494],db_even.mem_bank[2494]);
$fdisplay(file, "0x137E0,0x%h_0x%h", db_odd.mem_bank[2495],db_even.mem_bank[2495]);
$fdisplay(file, "0x13800,0x%h_0x%h", db_odd.mem_bank[2496],db_even.mem_bank[2496]);
$fdisplay(file, "0x13820,0x%h_0x%h", db_odd.mem_bank[2497],db_even.mem_bank[2497]);
$fdisplay(file, "0x13840,0x%h_0x%h", db_odd.mem_bank[2498],db_even.mem_bank[2498]);
$fdisplay(file, "0x13860,0x%h_0x%h", db_odd.mem_bank[2499],db_even.mem_bank[2499]);
$fdisplay(file, "0x13880,0x%h_0x%h", db_odd.mem_bank[2500],db_even.mem_bank[2500]);
$fdisplay(file, "0x138A0,0x%h_0x%h", db_odd.mem_bank[2501],db_even.mem_bank[2501]);
$fdisplay(file, "0x138C0,0x%h_0x%h", db_odd.mem_bank[2502],db_even.mem_bank[2502]);
$fdisplay(file, "0x138E0,0x%h_0x%h", db_odd.mem_bank[2503],db_even.mem_bank[2503]);
$fdisplay(file, "0x13900,0x%h_0x%h", db_odd.mem_bank[2504],db_even.mem_bank[2504]);
$fdisplay(file, "0x13920,0x%h_0x%h", db_odd.mem_bank[2505],db_even.mem_bank[2505]);
$fdisplay(file, "0x13940,0x%h_0x%h", db_odd.mem_bank[2506],db_even.mem_bank[2506]);
$fdisplay(file, "0x13960,0x%h_0x%h", db_odd.mem_bank[2507],db_even.mem_bank[2507]);
$fdisplay(file, "0x13980,0x%h_0x%h", db_odd.mem_bank[2508],db_even.mem_bank[2508]);
$fdisplay(file, "0x139A0,0x%h_0x%h", db_odd.mem_bank[2509],db_even.mem_bank[2509]);
$fdisplay(file, "0x139C0,0x%h_0x%h", db_odd.mem_bank[2510],db_even.mem_bank[2510]);
$fdisplay(file, "0x139E0,0x%h_0x%h", db_odd.mem_bank[2511],db_even.mem_bank[2511]);
$fdisplay(file, "0x13A00,0x%h_0x%h", db_odd.mem_bank[2512],db_even.mem_bank[2512]);
$fdisplay(file, "0x13A20,0x%h_0x%h", db_odd.mem_bank[2513],db_even.mem_bank[2513]);
$fdisplay(file, "0x13A40,0x%h_0x%h", db_odd.mem_bank[2514],db_even.mem_bank[2514]);
$fdisplay(file, "0x13A60,0x%h_0x%h", db_odd.mem_bank[2515],db_even.mem_bank[2515]);
$fdisplay(file, "0x13A80,0x%h_0x%h", db_odd.mem_bank[2516],db_even.mem_bank[2516]);
$fdisplay(file, "0x13AA0,0x%h_0x%h", db_odd.mem_bank[2517],db_even.mem_bank[2517]);
$fdisplay(file, "0x13AC0,0x%h_0x%h", db_odd.mem_bank[2518],db_even.mem_bank[2518]);
$fdisplay(file, "0x13AE0,0x%h_0x%h", db_odd.mem_bank[2519],db_even.mem_bank[2519]);
$fdisplay(file, "0x13B00,0x%h_0x%h", db_odd.mem_bank[2520],db_even.mem_bank[2520]);
$fdisplay(file, "0x13B20,0x%h_0x%h", db_odd.mem_bank[2521],db_even.mem_bank[2521]);
$fdisplay(file, "0x13B40,0x%h_0x%h", db_odd.mem_bank[2522],db_even.mem_bank[2522]);
$fdisplay(file, "0x13B60,0x%h_0x%h", db_odd.mem_bank[2523],db_even.mem_bank[2523]);
$fdisplay(file, "0x13B80,0x%h_0x%h", db_odd.mem_bank[2524],db_even.mem_bank[2524]);
$fdisplay(file, "0x13BA0,0x%h_0x%h", db_odd.mem_bank[2525],db_even.mem_bank[2525]);
$fdisplay(file, "0x13BC0,0x%h_0x%h", db_odd.mem_bank[2526],db_even.mem_bank[2526]);
$fdisplay(file, "0x13BE0,0x%h_0x%h", db_odd.mem_bank[2527],db_even.mem_bank[2527]);
$fdisplay(file, "0x13C00,0x%h_0x%h", db_odd.mem_bank[2528],db_even.mem_bank[2528]);
$fdisplay(file, "0x13C20,0x%h_0x%h", db_odd.mem_bank[2529],db_even.mem_bank[2529]);
$fdisplay(file, "0x13C40,0x%h_0x%h", db_odd.mem_bank[2530],db_even.mem_bank[2530]);
$fdisplay(file, "0x13C60,0x%h_0x%h", db_odd.mem_bank[2531],db_even.mem_bank[2531]);
$fdisplay(file, "0x13C80,0x%h_0x%h", db_odd.mem_bank[2532],db_even.mem_bank[2532]);
$fdisplay(file, "0x13CA0,0x%h_0x%h", db_odd.mem_bank[2533],db_even.mem_bank[2533]);
$fdisplay(file, "0x13CC0,0x%h_0x%h", db_odd.mem_bank[2534],db_even.mem_bank[2534]);
$fdisplay(file, "0x13CE0,0x%h_0x%h", db_odd.mem_bank[2535],db_even.mem_bank[2535]);
$fdisplay(file, "0x13D00,0x%h_0x%h", db_odd.mem_bank[2536],db_even.mem_bank[2536]);
$fdisplay(file, "0x13D20,0x%h_0x%h", db_odd.mem_bank[2537],db_even.mem_bank[2537]);
$fdisplay(file, "0x13D40,0x%h_0x%h", db_odd.mem_bank[2538],db_even.mem_bank[2538]);
$fdisplay(file, "0x13D60,0x%h_0x%h", db_odd.mem_bank[2539],db_even.mem_bank[2539]);
$fdisplay(file, "0x13D80,0x%h_0x%h", db_odd.mem_bank[2540],db_even.mem_bank[2540]);
$fdisplay(file, "0x13DA0,0x%h_0x%h", db_odd.mem_bank[2541],db_even.mem_bank[2541]);
$fdisplay(file, "0x13DC0,0x%h_0x%h", db_odd.mem_bank[2542],db_even.mem_bank[2542]);
$fdisplay(file, "0x13DE0,0x%h_0x%h", db_odd.mem_bank[2543],db_even.mem_bank[2543]);
$fdisplay(file, "0x13E00,0x%h_0x%h", db_odd.mem_bank[2544],db_even.mem_bank[2544]);
$fdisplay(file, "0x13E20,0x%h_0x%h", db_odd.mem_bank[2545],db_even.mem_bank[2545]);
$fdisplay(file, "0x13E40,0x%h_0x%h", db_odd.mem_bank[2546],db_even.mem_bank[2546]);
$fdisplay(file, "0x13E60,0x%h_0x%h", db_odd.mem_bank[2547],db_even.mem_bank[2547]);
$fdisplay(file, "0x13E80,0x%h_0x%h", db_odd.mem_bank[2548],db_even.mem_bank[2548]);
$fdisplay(file, "0x13EA0,0x%h_0x%h", db_odd.mem_bank[2549],db_even.mem_bank[2549]);
$fdisplay(file, "0x13EC0,0x%h_0x%h", db_odd.mem_bank[2550],db_even.mem_bank[2550]);
$fdisplay(file, "0x13EE0,0x%h_0x%h", db_odd.mem_bank[2551],db_even.mem_bank[2551]);
$fdisplay(file, "0x13F00,0x%h_0x%h", db_odd.mem_bank[2552],db_even.mem_bank[2552]);
$fdisplay(file, "0x13F20,0x%h_0x%h", db_odd.mem_bank[2553],db_even.mem_bank[2553]);
$fdisplay(file, "0x13F40,0x%h_0x%h", db_odd.mem_bank[2554],db_even.mem_bank[2554]);
$fdisplay(file, "0x13F60,0x%h_0x%h", db_odd.mem_bank[2555],db_even.mem_bank[2555]);
$fdisplay(file, "0x13F80,0x%h_0x%h", db_odd.mem_bank[2556],db_even.mem_bank[2556]);
$fdisplay(file, "0x13FA0,0x%h_0x%h", db_odd.mem_bank[2557],db_even.mem_bank[2557]);
$fdisplay(file, "0x13FC0,0x%h_0x%h", db_odd.mem_bank[2558],db_even.mem_bank[2558]);
$fdisplay(file, "0x13FE0,0x%h_0x%h", db_odd.mem_bank[2559],db_even.mem_bank[2559]);
$fdisplay(file, "0x14000,0x%h_0x%h", db_odd.mem_bank[2560],db_even.mem_bank[2560]);
$fdisplay(file, "0x14020,0x%h_0x%h", db_odd.mem_bank[2561],db_even.mem_bank[2561]);
$fdisplay(file, "0x14040,0x%h_0x%h", db_odd.mem_bank[2562],db_even.mem_bank[2562]);
$fdisplay(file, "0x14060,0x%h_0x%h", db_odd.mem_bank[2563],db_even.mem_bank[2563]);
$fdisplay(file, "0x14080,0x%h_0x%h", db_odd.mem_bank[2564],db_even.mem_bank[2564]);
$fdisplay(file, "0x140A0,0x%h_0x%h", db_odd.mem_bank[2565],db_even.mem_bank[2565]);
$fdisplay(file, "0x140C0,0x%h_0x%h", db_odd.mem_bank[2566],db_even.mem_bank[2566]);
$fdisplay(file, "0x140E0,0x%h_0x%h", db_odd.mem_bank[2567],db_even.mem_bank[2567]);
$fdisplay(file, "0x14100,0x%h_0x%h", db_odd.mem_bank[2568],db_even.mem_bank[2568]);
$fdisplay(file, "0x14120,0x%h_0x%h", db_odd.mem_bank[2569],db_even.mem_bank[2569]);
$fdisplay(file, "0x14140,0x%h_0x%h", db_odd.mem_bank[2570],db_even.mem_bank[2570]);
$fdisplay(file, "0x14160,0x%h_0x%h", db_odd.mem_bank[2571],db_even.mem_bank[2571]);
$fdisplay(file, "0x14180,0x%h_0x%h", db_odd.mem_bank[2572],db_even.mem_bank[2572]);
$fdisplay(file, "0x141A0,0x%h_0x%h", db_odd.mem_bank[2573],db_even.mem_bank[2573]);
$fdisplay(file, "0x141C0,0x%h_0x%h", db_odd.mem_bank[2574],db_even.mem_bank[2574]);
$fdisplay(file, "0x141E0,0x%h_0x%h", db_odd.mem_bank[2575],db_even.mem_bank[2575]);
$fdisplay(file, "0x14200,0x%h_0x%h", db_odd.mem_bank[2576],db_even.mem_bank[2576]);
$fdisplay(file, "0x14220,0x%h_0x%h", db_odd.mem_bank[2577],db_even.mem_bank[2577]);
$fdisplay(file, "0x14240,0x%h_0x%h", db_odd.mem_bank[2578],db_even.mem_bank[2578]);
$fdisplay(file, "0x14260,0x%h_0x%h", db_odd.mem_bank[2579],db_even.mem_bank[2579]);
$fdisplay(file, "0x14280,0x%h_0x%h", db_odd.mem_bank[2580],db_even.mem_bank[2580]);
$fdisplay(file, "0x142A0,0x%h_0x%h", db_odd.mem_bank[2581],db_even.mem_bank[2581]);
$fdisplay(file, "0x142C0,0x%h_0x%h", db_odd.mem_bank[2582],db_even.mem_bank[2582]);
$fdisplay(file, "0x142E0,0x%h_0x%h", db_odd.mem_bank[2583],db_even.mem_bank[2583]);
$fdisplay(file, "0x14300,0x%h_0x%h", db_odd.mem_bank[2584],db_even.mem_bank[2584]);
$fdisplay(file, "0x14320,0x%h_0x%h", db_odd.mem_bank[2585],db_even.mem_bank[2585]);
$fdisplay(file, "0x14340,0x%h_0x%h", db_odd.mem_bank[2586],db_even.mem_bank[2586]);
$fdisplay(file, "0x14360,0x%h_0x%h", db_odd.mem_bank[2587],db_even.mem_bank[2587]);
$fdisplay(file, "0x14380,0x%h_0x%h", db_odd.mem_bank[2588],db_even.mem_bank[2588]);
$fdisplay(file, "0x143A0,0x%h_0x%h", db_odd.mem_bank[2589],db_even.mem_bank[2589]);
$fdisplay(file, "0x143C0,0x%h_0x%h", db_odd.mem_bank[2590],db_even.mem_bank[2590]);
$fdisplay(file, "0x143E0,0x%h_0x%h", db_odd.mem_bank[2591],db_even.mem_bank[2591]);
$fdisplay(file, "0x14400,0x%h_0x%h", db_odd.mem_bank[2592],db_even.mem_bank[2592]);
$fdisplay(file, "0x14420,0x%h_0x%h", db_odd.mem_bank[2593],db_even.mem_bank[2593]);
$fdisplay(file, "0x14440,0x%h_0x%h", db_odd.mem_bank[2594],db_even.mem_bank[2594]);
$fdisplay(file, "0x14460,0x%h_0x%h", db_odd.mem_bank[2595],db_even.mem_bank[2595]);
$fdisplay(file, "0x14480,0x%h_0x%h", db_odd.mem_bank[2596],db_even.mem_bank[2596]);
$fdisplay(file, "0x144A0,0x%h_0x%h", db_odd.mem_bank[2597],db_even.mem_bank[2597]);
$fdisplay(file, "0x144C0,0x%h_0x%h", db_odd.mem_bank[2598],db_even.mem_bank[2598]);
$fdisplay(file, "0x144E0,0x%h_0x%h", db_odd.mem_bank[2599],db_even.mem_bank[2599]);
$fdisplay(file, "0x14500,0x%h_0x%h", db_odd.mem_bank[2600],db_even.mem_bank[2600]);
$fdisplay(file, "0x14520,0x%h_0x%h", db_odd.mem_bank[2601],db_even.mem_bank[2601]);
$fdisplay(file, "0x14540,0x%h_0x%h", db_odd.mem_bank[2602],db_even.mem_bank[2602]);
$fdisplay(file, "0x14560,0x%h_0x%h", db_odd.mem_bank[2603],db_even.mem_bank[2603]);
$fdisplay(file, "0x14580,0x%h_0x%h", db_odd.mem_bank[2604],db_even.mem_bank[2604]);
$fdisplay(file, "0x145A0,0x%h_0x%h", db_odd.mem_bank[2605],db_even.mem_bank[2605]);
$fdisplay(file, "0x145C0,0x%h_0x%h", db_odd.mem_bank[2606],db_even.mem_bank[2606]);
$fdisplay(file, "0x145E0,0x%h_0x%h", db_odd.mem_bank[2607],db_even.mem_bank[2607]);
$fdisplay(file, "0x14600,0x%h_0x%h", db_odd.mem_bank[2608],db_even.mem_bank[2608]);
$fdisplay(file, "0x14620,0x%h_0x%h", db_odd.mem_bank[2609],db_even.mem_bank[2609]);
$fdisplay(file, "0x14640,0x%h_0x%h", db_odd.mem_bank[2610],db_even.mem_bank[2610]);
$fdisplay(file, "0x14660,0x%h_0x%h", db_odd.mem_bank[2611],db_even.mem_bank[2611]);
$fdisplay(file, "0x14680,0x%h_0x%h", db_odd.mem_bank[2612],db_even.mem_bank[2612]);
$fdisplay(file, "0x146A0,0x%h_0x%h", db_odd.mem_bank[2613],db_even.mem_bank[2613]);
$fdisplay(file, "0x146C0,0x%h_0x%h", db_odd.mem_bank[2614],db_even.mem_bank[2614]);
$fdisplay(file, "0x146E0,0x%h_0x%h", db_odd.mem_bank[2615],db_even.mem_bank[2615]);
$fdisplay(file, "0x14700,0x%h_0x%h", db_odd.mem_bank[2616],db_even.mem_bank[2616]);
$fdisplay(file, "0x14720,0x%h_0x%h", db_odd.mem_bank[2617],db_even.mem_bank[2617]);
$fdisplay(file, "0x14740,0x%h_0x%h", db_odd.mem_bank[2618],db_even.mem_bank[2618]);
$fdisplay(file, "0x14760,0x%h_0x%h", db_odd.mem_bank[2619],db_even.mem_bank[2619]);
$fdisplay(file, "0x14780,0x%h_0x%h", db_odd.mem_bank[2620],db_even.mem_bank[2620]);
$fdisplay(file, "0x147A0,0x%h_0x%h", db_odd.mem_bank[2621],db_even.mem_bank[2621]);
$fdisplay(file, "0x147C0,0x%h_0x%h", db_odd.mem_bank[2622],db_even.mem_bank[2622]);
$fdisplay(file, "0x147E0,0x%h_0x%h", db_odd.mem_bank[2623],db_even.mem_bank[2623]);
$fdisplay(file, "0x14800,0x%h_0x%h", db_odd.mem_bank[2624],db_even.mem_bank[2624]);
$fdisplay(file, "0x14820,0x%h_0x%h", db_odd.mem_bank[2625],db_even.mem_bank[2625]);
$fdisplay(file, "0x14840,0x%h_0x%h", db_odd.mem_bank[2626],db_even.mem_bank[2626]);
$fdisplay(file, "0x14860,0x%h_0x%h", db_odd.mem_bank[2627],db_even.mem_bank[2627]);
$fdisplay(file, "0x14880,0x%h_0x%h", db_odd.mem_bank[2628],db_even.mem_bank[2628]);
$fdisplay(file, "0x148A0,0x%h_0x%h", db_odd.mem_bank[2629],db_even.mem_bank[2629]);
$fdisplay(file, "0x148C0,0x%h_0x%h", db_odd.mem_bank[2630],db_even.mem_bank[2630]);
$fdisplay(file, "0x148E0,0x%h_0x%h", db_odd.mem_bank[2631],db_even.mem_bank[2631]);
$fdisplay(file, "0x14900,0x%h_0x%h", db_odd.mem_bank[2632],db_even.mem_bank[2632]);
$fdisplay(file, "0x14920,0x%h_0x%h", db_odd.mem_bank[2633],db_even.mem_bank[2633]);
$fdisplay(file, "0x14940,0x%h_0x%h", db_odd.mem_bank[2634],db_even.mem_bank[2634]);
$fdisplay(file, "0x14960,0x%h_0x%h", db_odd.mem_bank[2635],db_even.mem_bank[2635]);
$fdisplay(file, "0x14980,0x%h_0x%h", db_odd.mem_bank[2636],db_even.mem_bank[2636]);
$fdisplay(file, "0x149A0,0x%h_0x%h", db_odd.mem_bank[2637],db_even.mem_bank[2637]);
$fdisplay(file, "0x149C0,0x%h_0x%h", db_odd.mem_bank[2638],db_even.mem_bank[2638]);
$fdisplay(file, "0x149E0,0x%h_0x%h", db_odd.mem_bank[2639],db_even.mem_bank[2639]);
$fdisplay(file, "0x14A00,0x%h_0x%h", db_odd.mem_bank[2640],db_even.mem_bank[2640]);
$fdisplay(file, "0x14A20,0x%h_0x%h", db_odd.mem_bank[2641],db_even.mem_bank[2641]);
$fdisplay(file, "0x14A40,0x%h_0x%h", db_odd.mem_bank[2642],db_even.mem_bank[2642]);
$fdisplay(file, "0x14A60,0x%h_0x%h", db_odd.mem_bank[2643],db_even.mem_bank[2643]);
$fdisplay(file, "0x14A80,0x%h_0x%h", db_odd.mem_bank[2644],db_even.mem_bank[2644]);
$fdisplay(file, "0x14AA0,0x%h_0x%h", db_odd.mem_bank[2645],db_even.mem_bank[2645]);
$fdisplay(file, "0x14AC0,0x%h_0x%h", db_odd.mem_bank[2646],db_even.mem_bank[2646]);
$fdisplay(file, "0x14AE0,0x%h_0x%h", db_odd.mem_bank[2647],db_even.mem_bank[2647]);
$fdisplay(file, "0x14B00,0x%h_0x%h", db_odd.mem_bank[2648],db_even.mem_bank[2648]);
$fdisplay(file, "0x14B20,0x%h_0x%h", db_odd.mem_bank[2649],db_even.mem_bank[2649]);
$fdisplay(file, "0x14B40,0x%h_0x%h", db_odd.mem_bank[2650],db_even.mem_bank[2650]);
$fdisplay(file, "0x14B60,0x%h_0x%h", db_odd.mem_bank[2651],db_even.mem_bank[2651]);
$fdisplay(file, "0x14B80,0x%h_0x%h", db_odd.mem_bank[2652],db_even.mem_bank[2652]);
$fdisplay(file, "0x14BA0,0x%h_0x%h", db_odd.mem_bank[2653],db_even.mem_bank[2653]);
$fdisplay(file, "0x14BC0,0x%h_0x%h", db_odd.mem_bank[2654],db_even.mem_bank[2654]);
$fdisplay(file, "0x14BE0,0x%h_0x%h", db_odd.mem_bank[2655],db_even.mem_bank[2655]);
$fdisplay(file, "0x14C00,0x%h_0x%h", db_odd.mem_bank[2656],db_even.mem_bank[2656]);
$fdisplay(file, "0x14C20,0x%h_0x%h", db_odd.mem_bank[2657],db_even.mem_bank[2657]);
$fdisplay(file, "0x14C40,0x%h_0x%h", db_odd.mem_bank[2658],db_even.mem_bank[2658]);
$fdisplay(file, "0x14C60,0x%h_0x%h", db_odd.mem_bank[2659],db_even.mem_bank[2659]);
$fdisplay(file, "0x14C80,0x%h_0x%h", db_odd.mem_bank[2660],db_even.mem_bank[2660]);
$fdisplay(file, "0x14CA0,0x%h_0x%h", db_odd.mem_bank[2661],db_even.mem_bank[2661]);
$fdisplay(file, "0x14CC0,0x%h_0x%h", db_odd.mem_bank[2662],db_even.mem_bank[2662]);
$fdisplay(file, "0x14CE0,0x%h_0x%h", db_odd.mem_bank[2663],db_even.mem_bank[2663]);
$fdisplay(file, "0x14D00,0x%h_0x%h", db_odd.mem_bank[2664],db_even.mem_bank[2664]);
$fdisplay(file, "0x14D20,0x%h_0x%h", db_odd.mem_bank[2665],db_even.mem_bank[2665]);
$fdisplay(file, "0x14D40,0x%h_0x%h", db_odd.mem_bank[2666],db_even.mem_bank[2666]);
$fdisplay(file, "0x14D60,0x%h_0x%h", db_odd.mem_bank[2667],db_even.mem_bank[2667]);
$fdisplay(file, "0x14D80,0x%h_0x%h", db_odd.mem_bank[2668],db_even.mem_bank[2668]);
$fdisplay(file, "0x14DA0,0x%h_0x%h", db_odd.mem_bank[2669],db_even.mem_bank[2669]);
$fdisplay(file, "0x14DC0,0x%h_0x%h", db_odd.mem_bank[2670],db_even.mem_bank[2670]);
$fdisplay(file, "0x14DE0,0x%h_0x%h", db_odd.mem_bank[2671],db_even.mem_bank[2671]);
$fdisplay(file, "0x14E00,0x%h_0x%h", db_odd.mem_bank[2672],db_even.mem_bank[2672]);
$fdisplay(file, "0x14E20,0x%h_0x%h", db_odd.mem_bank[2673],db_even.mem_bank[2673]);
$fdisplay(file, "0x14E40,0x%h_0x%h", db_odd.mem_bank[2674],db_even.mem_bank[2674]);
$fdisplay(file, "0x14E60,0x%h_0x%h", db_odd.mem_bank[2675],db_even.mem_bank[2675]);
$fdisplay(file, "0x14E80,0x%h_0x%h", db_odd.mem_bank[2676],db_even.mem_bank[2676]);
$fdisplay(file, "0x14EA0,0x%h_0x%h", db_odd.mem_bank[2677],db_even.mem_bank[2677]);
$fdisplay(file, "0x14EC0,0x%h_0x%h", db_odd.mem_bank[2678],db_even.mem_bank[2678]);
$fdisplay(file, "0x14EE0,0x%h_0x%h", db_odd.mem_bank[2679],db_even.mem_bank[2679]);
$fdisplay(file, "0x14F00,0x%h_0x%h", db_odd.mem_bank[2680],db_even.mem_bank[2680]);
$fdisplay(file, "0x14F20,0x%h_0x%h", db_odd.mem_bank[2681],db_even.mem_bank[2681]);
$fdisplay(file, "0x14F40,0x%h_0x%h", db_odd.mem_bank[2682],db_even.mem_bank[2682]);
$fdisplay(file, "0x14F60,0x%h_0x%h", db_odd.mem_bank[2683],db_even.mem_bank[2683]);
$fdisplay(file, "0x14F80,0x%h_0x%h", db_odd.mem_bank[2684],db_even.mem_bank[2684]);
$fdisplay(file, "0x14FA0,0x%h_0x%h", db_odd.mem_bank[2685],db_even.mem_bank[2685]);
$fdisplay(file, "0x14FC0,0x%h_0x%h", db_odd.mem_bank[2686],db_even.mem_bank[2686]);
$fdisplay(file, "0x14FE0,0x%h_0x%h", db_odd.mem_bank[2687],db_even.mem_bank[2687]);
$fdisplay(file, "0x15000,0x%h_0x%h", db_odd.mem_bank[2688],db_even.mem_bank[2688]);
$fdisplay(file, "0x15020,0x%h_0x%h", db_odd.mem_bank[2689],db_even.mem_bank[2689]);
$fdisplay(file, "0x15040,0x%h_0x%h", db_odd.mem_bank[2690],db_even.mem_bank[2690]);
$fdisplay(file, "0x15060,0x%h_0x%h", db_odd.mem_bank[2691],db_even.mem_bank[2691]);
$fdisplay(file, "0x15080,0x%h_0x%h", db_odd.mem_bank[2692],db_even.mem_bank[2692]);
$fdisplay(file, "0x150A0,0x%h_0x%h", db_odd.mem_bank[2693],db_even.mem_bank[2693]);
$fdisplay(file, "0x150C0,0x%h_0x%h", db_odd.mem_bank[2694],db_even.mem_bank[2694]);
$fdisplay(file, "0x150E0,0x%h_0x%h", db_odd.mem_bank[2695],db_even.mem_bank[2695]);
$fdisplay(file, "0x15100,0x%h_0x%h", db_odd.mem_bank[2696],db_even.mem_bank[2696]);
$fdisplay(file, "0x15120,0x%h_0x%h", db_odd.mem_bank[2697],db_even.mem_bank[2697]);
$fdisplay(file, "0x15140,0x%h_0x%h", db_odd.mem_bank[2698],db_even.mem_bank[2698]);
$fdisplay(file, "0x15160,0x%h_0x%h", db_odd.mem_bank[2699],db_even.mem_bank[2699]);
$fdisplay(file, "0x15180,0x%h_0x%h", db_odd.mem_bank[2700],db_even.mem_bank[2700]);
$fdisplay(file, "0x151A0,0x%h_0x%h", db_odd.mem_bank[2701],db_even.mem_bank[2701]);
$fdisplay(file, "0x151C0,0x%h_0x%h", db_odd.mem_bank[2702],db_even.mem_bank[2702]);
$fdisplay(file, "0x151E0,0x%h_0x%h", db_odd.mem_bank[2703],db_even.mem_bank[2703]);
$fdisplay(file, "0x15200,0x%h_0x%h", db_odd.mem_bank[2704],db_even.mem_bank[2704]);
$fdisplay(file, "0x15220,0x%h_0x%h", db_odd.mem_bank[2705],db_even.mem_bank[2705]);
$fdisplay(file, "0x15240,0x%h_0x%h", db_odd.mem_bank[2706],db_even.mem_bank[2706]);
$fdisplay(file, "0x15260,0x%h_0x%h", db_odd.mem_bank[2707],db_even.mem_bank[2707]);
$fdisplay(file, "0x15280,0x%h_0x%h", db_odd.mem_bank[2708],db_even.mem_bank[2708]);
$fdisplay(file, "0x152A0,0x%h_0x%h", db_odd.mem_bank[2709],db_even.mem_bank[2709]);
$fdisplay(file, "0x152C0,0x%h_0x%h", db_odd.mem_bank[2710],db_even.mem_bank[2710]);
$fdisplay(file, "0x152E0,0x%h_0x%h", db_odd.mem_bank[2711],db_even.mem_bank[2711]);
$fdisplay(file, "0x15300,0x%h_0x%h", db_odd.mem_bank[2712],db_even.mem_bank[2712]);
$fdisplay(file, "0x15320,0x%h_0x%h", db_odd.mem_bank[2713],db_even.mem_bank[2713]);
$fdisplay(file, "0x15340,0x%h_0x%h", db_odd.mem_bank[2714],db_even.mem_bank[2714]);
$fdisplay(file, "0x15360,0x%h_0x%h", db_odd.mem_bank[2715],db_even.mem_bank[2715]);
$fdisplay(file, "0x15380,0x%h_0x%h", db_odd.mem_bank[2716],db_even.mem_bank[2716]);
$fdisplay(file, "0x153A0,0x%h_0x%h", db_odd.mem_bank[2717],db_even.mem_bank[2717]);
$fdisplay(file, "0x153C0,0x%h_0x%h", db_odd.mem_bank[2718],db_even.mem_bank[2718]);
$fdisplay(file, "0x153E0,0x%h_0x%h", db_odd.mem_bank[2719],db_even.mem_bank[2719]);
$fdisplay(file, "0x15400,0x%h_0x%h", db_odd.mem_bank[2720],db_even.mem_bank[2720]);
$fdisplay(file, "0x15420,0x%h_0x%h", db_odd.mem_bank[2721],db_even.mem_bank[2721]);
$fdisplay(file, "0x15440,0x%h_0x%h", db_odd.mem_bank[2722],db_even.mem_bank[2722]);
$fdisplay(file, "0x15460,0x%h_0x%h", db_odd.mem_bank[2723],db_even.mem_bank[2723]);
$fdisplay(file, "0x15480,0x%h_0x%h", db_odd.mem_bank[2724],db_even.mem_bank[2724]);
$fdisplay(file, "0x154A0,0x%h_0x%h", db_odd.mem_bank[2725],db_even.mem_bank[2725]);
$fdisplay(file, "0x154C0,0x%h_0x%h", db_odd.mem_bank[2726],db_even.mem_bank[2726]);
$fdisplay(file, "0x154E0,0x%h_0x%h", db_odd.mem_bank[2727],db_even.mem_bank[2727]);
$fdisplay(file, "0x15500,0x%h_0x%h", db_odd.mem_bank[2728],db_even.mem_bank[2728]);
$fdisplay(file, "0x15520,0x%h_0x%h", db_odd.mem_bank[2729],db_even.mem_bank[2729]);
$fdisplay(file, "0x15540,0x%h_0x%h", db_odd.mem_bank[2730],db_even.mem_bank[2730]);
$fdisplay(file, "0x15560,0x%h_0x%h", db_odd.mem_bank[2731],db_even.mem_bank[2731]);
$fdisplay(file, "0x15580,0x%h_0x%h", db_odd.mem_bank[2732],db_even.mem_bank[2732]);
$fdisplay(file, "0x155A0,0x%h_0x%h", db_odd.mem_bank[2733],db_even.mem_bank[2733]);
$fdisplay(file, "0x155C0,0x%h_0x%h", db_odd.mem_bank[2734],db_even.mem_bank[2734]);
$fdisplay(file, "0x155E0,0x%h_0x%h", db_odd.mem_bank[2735],db_even.mem_bank[2735]);
$fdisplay(file, "0x15600,0x%h_0x%h", db_odd.mem_bank[2736],db_even.mem_bank[2736]);
$fdisplay(file, "0x15620,0x%h_0x%h", db_odd.mem_bank[2737],db_even.mem_bank[2737]);
$fdisplay(file, "0x15640,0x%h_0x%h", db_odd.mem_bank[2738],db_even.mem_bank[2738]);
$fdisplay(file, "0x15660,0x%h_0x%h", db_odd.mem_bank[2739],db_even.mem_bank[2739]);
$fdisplay(file, "0x15680,0x%h_0x%h", db_odd.mem_bank[2740],db_even.mem_bank[2740]);
$fdisplay(file, "0x156A0,0x%h_0x%h", db_odd.mem_bank[2741],db_even.mem_bank[2741]);
$fdisplay(file, "0x156C0,0x%h_0x%h", db_odd.mem_bank[2742],db_even.mem_bank[2742]);
$fdisplay(file, "0x156E0,0x%h_0x%h", db_odd.mem_bank[2743],db_even.mem_bank[2743]);
$fdisplay(file, "0x15700,0x%h_0x%h", db_odd.mem_bank[2744],db_even.mem_bank[2744]);
$fdisplay(file, "0x15720,0x%h_0x%h", db_odd.mem_bank[2745],db_even.mem_bank[2745]);
$fdisplay(file, "0x15740,0x%h_0x%h", db_odd.mem_bank[2746],db_even.mem_bank[2746]);
$fdisplay(file, "0x15760,0x%h_0x%h", db_odd.mem_bank[2747],db_even.mem_bank[2747]);
$fdisplay(file, "0x15780,0x%h_0x%h", db_odd.mem_bank[2748],db_even.mem_bank[2748]);
$fdisplay(file, "0x157A0,0x%h_0x%h", db_odd.mem_bank[2749],db_even.mem_bank[2749]);
$fdisplay(file, "0x157C0,0x%h_0x%h", db_odd.mem_bank[2750],db_even.mem_bank[2750]);
$fdisplay(file, "0x157E0,0x%h_0x%h", db_odd.mem_bank[2751],db_even.mem_bank[2751]);
$fdisplay(file, "0x15800,0x%h_0x%h", db_odd.mem_bank[2752],db_even.mem_bank[2752]);
$fdisplay(file, "0x15820,0x%h_0x%h", db_odd.mem_bank[2753],db_even.mem_bank[2753]);
$fdisplay(file, "0x15840,0x%h_0x%h", db_odd.mem_bank[2754],db_even.mem_bank[2754]);
$fdisplay(file, "0x15860,0x%h_0x%h", db_odd.mem_bank[2755],db_even.mem_bank[2755]);
$fdisplay(file, "0x15880,0x%h_0x%h", db_odd.mem_bank[2756],db_even.mem_bank[2756]);
$fdisplay(file, "0x158A0,0x%h_0x%h", db_odd.mem_bank[2757],db_even.mem_bank[2757]);
$fdisplay(file, "0x158C0,0x%h_0x%h", db_odd.mem_bank[2758],db_even.mem_bank[2758]);
$fdisplay(file, "0x158E0,0x%h_0x%h", db_odd.mem_bank[2759],db_even.mem_bank[2759]);
$fdisplay(file, "0x15900,0x%h_0x%h", db_odd.mem_bank[2760],db_even.mem_bank[2760]);
$fdisplay(file, "0x15920,0x%h_0x%h", db_odd.mem_bank[2761],db_even.mem_bank[2761]);
$fdisplay(file, "0x15940,0x%h_0x%h", db_odd.mem_bank[2762],db_even.mem_bank[2762]);
$fdisplay(file, "0x15960,0x%h_0x%h", db_odd.mem_bank[2763],db_even.mem_bank[2763]);
$fdisplay(file, "0x15980,0x%h_0x%h", db_odd.mem_bank[2764],db_even.mem_bank[2764]);
$fdisplay(file, "0x159A0,0x%h_0x%h", db_odd.mem_bank[2765],db_even.mem_bank[2765]);
$fdisplay(file, "0x159C0,0x%h_0x%h", db_odd.mem_bank[2766],db_even.mem_bank[2766]);
$fdisplay(file, "0x159E0,0x%h_0x%h", db_odd.mem_bank[2767],db_even.mem_bank[2767]);
$fdisplay(file, "0x15A00,0x%h_0x%h", db_odd.mem_bank[2768],db_even.mem_bank[2768]);
$fdisplay(file, "0x15A20,0x%h_0x%h", db_odd.mem_bank[2769],db_even.mem_bank[2769]);
$fdisplay(file, "0x15A40,0x%h_0x%h", db_odd.mem_bank[2770],db_even.mem_bank[2770]);
$fdisplay(file, "0x15A60,0x%h_0x%h", db_odd.mem_bank[2771],db_even.mem_bank[2771]);
$fdisplay(file, "0x15A80,0x%h_0x%h", db_odd.mem_bank[2772],db_even.mem_bank[2772]);
$fdisplay(file, "0x15AA0,0x%h_0x%h", db_odd.mem_bank[2773],db_even.mem_bank[2773]);
$fdisplay(file, "0x15AC0,0x%h_0x%h", db_odd.mem_bank[2774],db_even.mem_bank[2774]);
$fdisplay(file, "0x15AE0,0x%h_0x%h", db_odd.mem_bank[2775],db_even.mem_bank[2775]);
$fdisplay(file, "0x15B00,0x%h_0x%h", db_odd.mem_bank[2776],db_even.mem_bank[2776]);
$fdisplay(file, "0x15B20,0x%h_0x%h", db_odd.mem_bank[2777],db_even.mem_bank[2777]);
$fdisplay(file, "0x15B40,0x%h_0x%h", db_odd.mem_bank[2778],db_even.mem_bank[2778]);
$fdisplay(file, "0x15B60,0x%h_0x%h", db_odd.mem_bank[2779],db_even.mem_bank[2779]);
$fdisplay(file, "0x15B80,0x%h_0x%h", db_odd.mem_bank[2780],db_even.mem_bank[2780]);
$fdisplay(file, "0x15BA0,0x%h_0x%h", db_odd.mem_bank[2781],db_even.mem_bank[2781]);
$fdisplay(file, "0x15BC0,0x%h_0x%h", db_odd.mem_bank[2782],db_even.mem_bank[2782]);
$fdisplay(file, "0x15BE0,0x%h_0x%h", db_odd.mem_bank[2783],db_even.mem_bank[2783]);
$fdisplay(file, "0x15C00,0x%h_0x%h", db_odd.mem_bank[2784],db_even.mem_bank[2784]);
$fdisplay(file, "0x15C20,0x%h_0x%h", db_odd.mem_bank[2785],db_even.mem_bank[2785]);
$fdisplay(file, "0x15C40,0x%h_0x%h", db_odd.mem_bank[2786],db_even.mem_bank[2786]);
$fdisplay(file, "0x15C60,0x%h_0x%h", db_odd.mem_bank[2787],db_even.mem_bank[2787]);
$fdisplay(file, "0x15C80,0x%h_0x%h", db_odd.mem_bank[2788],db_even.mem_bank[2788]);
$fdisplay(file, "0x15CA0,0x%h_0x%h", db_odd.mem_bank[2789],db_even.mem_bank[2789]);
$fdisplay(file, "0x15CC0,0x%h_0x%h", db_odd.mem_bank[2790],db_even.mem_bank[2790]);
$fdisplay(file, "0x15CE0,0x%h_0x%h", db_odd.mem_bank[2791],db_even.mem_bank[2791]);
$fdisplay(file, "0x15D00,0x%h_0x%h", db_odd.mem_bank[2792],db_even.mem_bank[2792]);
$fdisplay(file, "0x15D20,0x%h_0x%h", db_odd.mem_bank[2793],db_even.mem_bank[2793]);
$fdisplay(file, "0x15D40,0x%h_0x%h", db_odd.mem_bank[2794],db_even.mem_bank[2794]);
$fdisplay(file, "0x15D60,0x%h_0x%h", db_odd.mem_bank[2795],db_even.mem_bank[2795]);
$fdisplay(file, "0x15D80,0x%h_0x%h", db_odd.mem_bank[2796],db_even.mem_bank[2796]);
$fdisplay(file, "0x15DA0,0x%h_0x%h", db_odd.mem_bank[2797],db_even.mem_bank[2797]);
$fdisplay(file, "0x15DC0,0x%h_0x%h", db_odd.mem_bank[2798],db_even.mem_bank[2798]);
$fdisplay(file, "0x15DE0,0x%h_0x%h", db_odd.mem_bank[2799],db_even.mem_bank[2799]);
$fdisplay(file, "0x15E00,0x%h_0x%h", db_odd.mem_bank[2800],db_even.mem_bank[2800]);
$fdisplay(file, "0x15E20,0x%h_0x%h", db_odd.mem_bank[2801],db_even.mem_bank[2801]);
$fdisplay(file, "0x15E40,0x%h_0x%h", db_odd.mem_bank[2802],db_even.mem_bank[2802]);
$fdisplay(file, "0x15E60,0x%h_0x%h", db_odd.mem_bank[2803],db_even.mem_bank[2803]);
$fdisplay(file, "0x15E80,0x%h_0x%h", db_odd.mem_bank[2804],db_even.mem_bank[2804]);
$fdisplay(file, "0x15EA0,0x%h_0x%h", db_odd.mem_bank[2805],db_even.mem_bank[2805]);
$fdisplay(file, "0x15EC0,0x%h_0x%h", db_odd.mem_bank[2806],db_even.mem_bank[2806]);
$fdisplay(file, "0x15EE0,0x%h_0x%h", db_odd.mem_bank[2807],db_even.mem_bank[2807]);
$fdisplay(file, "0x15F00,0x%h_0x%h", db_odd.mem_bank[2808],db_even.mem_bank[2808]);
$fdisplay(file, "0x15F20,0x%h_0x%h", db_odd.mem_bank[2809],db_even.mem_bank[2809]);
$fdisplay(file, "0x15F40,0x%h_0x%h", db_odd.mem_bank[2810],db_even.mem_bank[2810]);
$fdisplay(file, "0x15F60,0x%h_0x%h", db_odd.mem_bank[2811],db_even.mem_bank[2811]);
$fdisplay(file, "0x15F80,0x%h_0x%h", db_odd.mem_bank[2812],db_even.mem_bank[2812]);
$fdisplay(file, "0x15FA0,0x%h_0x%h", db_odd.mem_bank[2813],db_even.mem_bank[2813]);
$fdisplay(file, "0x15FC0,0x%h_0x%h", db_odd.mem_bank[2814],db_even.mem_bank[2814]);
$fdisplay(file, "0x15FE0,0x%h_0x%h", db_odd.mem_bank[2815],db_even.mem_bank[2815]);
$fdisplay(file, "0x16000,0x%h_0x%h", db_odd.mem_bank[2816],db_even.mem_bank[2816]);
$fdisplay(file, "0x16020,0x%h_0x%h", db_odd.mem_bank[2817],db_even.mem_bank[2817]);
$fdisplay(file, "0x16040,0x%h_0x%h", db_odd.mem_bank[2818],db_even.mem_bank[2818]);
$fdisplay(file, "0x16060,0x%h_0x%h", db_odd.mem_bank[2819],db_even.mem_bank[2819]);
$fdisplay(file, "0x16080,0x%h_0x%h", db_odd.mem_bank[2820],db_even.mem_bank[2820]);
$fdisplay(file, "0x160A0,0x%h_0x%h", db_odd.mem_bank[2821],db_even.mem_bank[2821]);
$fdisplay(file, "0x160C0,0x%h_0x%h", db_odd.mem_bank[2822],db_even.mem_bank[2822]);
$fdisplay(file, "0x160E0,0x%h_0x%h", db_odd.mem_bank[2823],db_even.mem_bank[2823]);
$fdisplay(file, "0x16100,0x%h_0x%h", db_odd.mem_bank[2824],db_even.mem_bank[2824]);
$fdisplay(file, "0x16120,0x%h_0x%h", db_odd.mem_bank[2825],db_even.mem_bank[2825]);
$fdisplay(file, "0x16140,0x%h_0x%h", db_odd.mem_bank[2826],db_even.mem_bank[2826]);
$fdisplay(file, "0x16160,0x%h_0x%h", db_odd.mem_bank[2827],db_even.mem_bank[2827]);
$fdisplay(file, "0x16180,0x%h_0x%h", db_odd.mem_bank[2828],db_even.mem_bank[2828]);
$fdisplay(file, "0x161A0,0x%h_0x%h", db_odd.mem_bank[2829],db_even.mem_bank[2829]);
$fdisplay(file, "0x161C0,0x%h_0x%h", db_odd.mem_bank[2830],db_even.mem_bank[2830]);
$fdisplay(file, "0x161E0,0x%h_0x%h", db_odd.mem_bank[2831],db_even.mem_bank[2831]);
$fdisplay(file, "0x16200,0x%h_0x%h", db_odd.mem_bank[2832],db_even.mem_bank[2832]);
$fdisplay(file, "0x16220,0x%h_0x%h", db_odd.mem_bank[2833],db_even.mem_bank[2833]);
$fdisplay(file, "0x16240,0x%h_0x%h", db_odd.mem_bank[2834],db_even.mem_bank[2834]);
$fdisplay(file, "0x16260,0x%h_0x%h", db_odd.mem_bank[2835],db_even.mem_bank[2835]);
$fdisplay(file, "0x16280,0x%h_0x%h", db_odd.mem_bank[2836],db_even.mem_bank[2836]);
$fdisplay(file, "0x162A0,0x%h_0x%h", db_odd.mem_bank[2837],db_even.mem_bank[2837]);
$fdisplay(file, "0x162C0,0x%h_0x%h", db_odd.mem_bank[2838],db_even.mem_bank[2838]);
$fdisplay(file, "0x162E0,0x%h_0x%h", db_odd.mem_bank[2839],db_even.mem_bank[2839]);
$fdisplay(file, "0x16300,0x%h_0x%h", db_odd.mem_bank[2840],db_even.mem_bank[2840]);
$fdisplay(file, "0x16320,0x%h_0x%h", db_odd.mem_bank[2841],db_even.mem_bank[2841]);
$fdisplay(file, "0x16340,0x%h_0x%h", db_odd.mem_bank[2842],db_even.mem_bank[2842]);
$fdisplay(file, "0x16360,0x%h_0x%h", db_odd.mem_bank[2843],db_even.mem_bank[2843]);
$fdisplay(file, "0x16380,0x%h_0x%h", db_odd.mem_bank[2844],db_even.mem_bank[2844]);
$fdisplay(file, "0x163A0,0x%h_0x%h", db_odd.mem_bank[2845],db_even.mem_bank[2845]);
$fdisplay(file, "0x163C0,0x%h_0x%h", db_odd.mem_bank[2846],db_even.mem_bank[2846]);
$fdisplay(file, "0x163E0,0x%h_0x%h", db_odd.mem_bank[2847],db_even.mem_bank[2847]);
$fdisplay(file, "0x16400,0x%h_0x%h", db_odd.mem_bank[2848],db_even.mem_bank[2848]);
$fdisplay(file, "0x16420,0x%h_0x%h", db_odd.mem_bank[2849],db_even.mem_bank[2849]);
$fdisplay(file, "0x16440,0x%h_0x%h", db_odd.mem_bank[2850],db_even.mem_bank[2850]);
$fdisplay(file, "0x16460,0x%h_0x%h", db_odd.mem_bank[2851],db_even.mem_bank[2851]);
$fdisplay(file, "0x16480,0x%h_0x%h", db_odd.mem_bank[2852],db_even.mem_bank[2852]);
$fdisplay(file, "0x164A0,0x%h_0x%h", db_odd.mem_bank[2853],db_even.mem_bank[2853]);
$fdisplay(file, "0x164C0,0x%h_0x%h", db_odd.mem_bank[2854],db_even.mem_bank[2854]);
$fdisplay(file, "0x164E0,0x%h_0x%h", db_odd.mem_bank[2855],db_even.mem_bank[2855]);
$fdisplay(file, "0x16500,0x%h_0x%h", db_odd.mem_bank[2856],db_even.mem_bank[2856]);
$fdisplay(file, "0x16520,0x%h_0x%h", db_odd.mem_bank[2857],db_even.mem_bank[2857]);
$fdisplay(file, "0x16540,0x%h_0x%h", db_odd.mem_bank[2858],db_even.mem_bank[2858]);
$fdisplay(file, "0x16560,0x%h_0x%h", db_odd.mem_bank[2859],db_even.mem_bank[2859]);
$fdisplay(file, "0x16580,0x%h_0x%h", db_odd.mem_bank[2860],db_even.mem_bank[2860]);
$fdisplay(file, "0x165A0,0x%h_0x%h", db_odd.mem_bank[2861],db_even.mem_bank[2861]);
$fdisplay(file, "0x165C0,0x%h_0x%h", db_odd.mem_bank[2862],db_even.mem_bank[2862]);
$fdisplay(file, "0x165E0,0x%h_0x%h", db_odd.mem_bank[2863],db_even.mem_bank[2863]);
$fdisplay(file, "0x16600,0x%h_0x%h", db_odd.mem_bank[2864],db_even.mem_bank[2864]);
$fdisplay(file, "0x16620,0x%h_0x%h", db_odd.mem_bank[2865],db_even.mem_bank[2865]);
$fdisplay(file, "0x16640,0x%h_0x%h", db_odd.mem_bank[2866],db_even.mem_bank[2866]);
$fdisplay(file, "0x16660,0x%h_0x%h", db_odd.mem_bank[2867],db_even.mem_bank[2867]);
$fdisplay(file, "0x16680,0x%h_0x%h", db_odd.mem_bank[2868],db_even.mem_bank[2868]);
$fdisplay(file, "0x166A0,0x%h_0x%h", db_odd.mem_bank[2869],db_even.mem_bank[2869]);
$fdisplay(file, "0x166C0,0x%h_0x%h", db_odd.mem_bank[2870],db_even.mem_bank[2870]);
$fdisplay(file, "0x166E0,0x%h_0x%h", db_odd.mem_bank[2871],db_even.mem_bank[2871]);
$fdisplay(file, "0x16700,0x%h_0x%h", db_odd.mem_bank[2872],db_even.mem_bank[2872]);
$fdisplay(file, "0x16720,0x%h_0x%h", db_odd.mem_bank[2873],db_even.mem_bank[2873]);
$fdisplay(file, "0x16740,0x%h_0x%h", db_odd.mem_bank[2874],db_even.mem_bank[2874]);
$fdisplay(file, "0x16760,0x%h_0x%h", db_odd.mem_bank[2875],db_even.mem_bank[2875]);
$fdisplay(file, "0x16780,0x%h_0x%h", db_odd.mem_bank[2876],db_even.mem_bank[2876]);
$fdisplay(file, "0x167A0,0x%h_0x%h", db_odd.mem_bank[2877],db_even.mem_bank[2877]);
$fdisplay(file, "0x167C0,0x%h_0x%h", db_odd.mem_bank[2878],db_even.mem_bank[2878]);
$fdisplay(file, "0x167E0,0x%h_0x%h", db_odd.mem_bank[2879],db_even.mem_bank[2879]);
$fdisplay(file, "0x16800,0x%h_0x%h", db_odd.mem_bank[2880],db_even.mem_bank[2880]);
$fdisplay(file, "0x16820,0x%h_0x%h", db_odd.mem_bank[2881],db_even.mem_bank[2881]);
$fdisplay(file, "0x16840,0x%h_0x%h", db_odd.mem_bank[2882],db_even.mem_bank[2882]);
$fdisplay(file, "0x16860,0x%h_0x%h", db_odd.mem_bank[2883],db_even.mem_bank[2883]);
$fdisplay(file, "0x16880,0x%h_0x%h", db_odd.mem_bank[2884],db_even.mem_bank[2884]);
$fdisplay(file, "0x168A0,0x%h_0x%h", db_odd.mem_bank[2885],db_even.mem_bank[2885]);
$fdisplay(file, "0x168C0,0x%h_0x%h", db_odd.mem_bank[2886],db_even.mem_bank[2886]);
$fdisplay(file, "0x168E0,0x%h_0x%h", db_odd.mem_bank[2887],db_even.mem_bank[2887]);
$fdisplay(file, "0x16900,0x%h_0x%h", db_odd.mem_bank[2888],db_even.mem_bank[2888]);
$fdisplay(file, "0x16920,0x%h_0x%h", db_odd.mem_bank[2889],db_even.mem_bank[2889]);
$fdisplay(file, "0x16940,0x%h_0x%h", db_odd.mem_bank[2890],db_even.mem_bank[2890]);
$fdisplay(file, "0x16960,0x%h_0x%h", db_odd.mem_bank[2891],db_even.mem_bank[2891]);
$fdisplay(file, "0x16980,0x%h_0x%h", db_odd.mem_bank[2892],db_even.mem_bank[2892]);
$fdisplay(file, "0x169A0,0x%h_0x%h", db_odd.mem_bank[2893],db_even.mem_bank[2893]);
$fdisplay(file, "0x169C0,0x%h_0x%h", db_odd.mem_bank[2894],db_even.mem_bank[2894]);
$fdisplay(file, "0x169E0,0x%h_0x%h", db_odd.mem_bank[2895],db_even.mem_bank[2895]);
$fdisplay(file, "0x16A00,0x%h_0x%h", db_odd.mem_bank[2896],db_even.mem_bank[2896]);
$fdisplay(file, "0x16A20,0x%h_0x%h", db_odd.mem_bank[2897],db_even.mem_bank[2897]);
$fdisplay(file, "0x16A40,0x%h_0x%h", db_odd.mem_bank[2898],db_even.mem_bank[2898]);
$fdisplay(file, "0x16A60,0x%h_0x%h", db_odd.mem_bank[2899],db_even.mem_bank[2899]);
$fdisplay(file, "0x16A80,0x%h_0x%h", db_odd.mem_bank[2900],db_even.mem_bank[2900]);
$fdisplay(file, "0x16AA0,0x%h_0x%h", db_odd.mem_bank[2901],db_even.mem_bank[2901]);
$fdisplay(file, "0x16AC0,0x%h_0x%h", db_odd.mem_bank[2902],db_even.mem_bank[2902]);
$fdisplay(file, "0x16AE0,0x%h_0x%h", db_odd.mem_bank[2903],db_even.mem_bank[2903]);
$fdisplay(file, "0x16B00,0x%h_0x%h", db_odd.mem_bank[2904],db_even.mem_bank[2904]);
$fdisplay(file, "0x16B20,0x%h_0x%h", db_odd.mem_bank[2905],db_even.mem_bank[2905]);
$fdisplay(file, "0x16B40,0x%h_0x%h", db_odd.mem_bank[2906],db_even.mem_bank[2906]);
$fdisplay(file, "0x16B60,0x%h_0x%h", db_odd.mem_bank[2907],db_even.mem_bank[2907]);
$fdisplay(file, "0x16B80,0x%h_0x%h", db_odd.mem_bank[2908],db_even.mem_bank[2908]);
$fdisplay(file, "0x16BA0,0x%h_0x%h", db_odd.mem_bank[2909],db_even.mem_bank[2909]);
$fdisplay(file, "0x16BC0,0x%h_0x%h", db_odd.mem_bank[2910],db_even.mem_bank[2910]);
$fdisplay(file, "0x16BE0,0x%h_0x%h", db_odd.mem_bank[2911],db_even.mem_bank[2911]);
$fdisplay(file, "0x16C00,0x%h_0x%h", db_odd.mem_bank[2912],db_even.mem_bank[2912]);
$fdisplay(file, "0x16C20,0x%h_0x%h", db_odd.mem_bank[2913],db_even.mem_bank[2913]);
$fdisplay(file, "0x16C40,0x%h_0x%h", db_odd.mem_bank[2914],db_even.mem_bank[2914]);
$fdisplay(file, "0x16C60,0x%h_0x%h", db_odd.mem_bank[2915],db_even.mem_bank[2915]);
$fdisplay(file, "0x16C80,0x%h_0x%h", db_odd.mem_bank[2916],db_even.mem_bank[2916]);
$fdisplay(file, "0x16CA0,0x%h_0x%h", db_odd.mem_bank[2917],db_even.mem_bank[2917]);
$fdisplay(file, "0x16CC0,0x%h_0x%h", db_odd.mem_bank[2918],db_even.mem_bank[2918]);
$fdisplay(file, "0x16CE0,0x%h_0x%h", db_odd.mem_bank[2919],db_even.mem_bank[2919]);
$fdisplay(file, "0x16D00,0x%h_0x%h", db_odd.mem_bank[2920],db_even.mem_bank[2920]);
$fdisplay(file, "0x16D20,0x%h_0x%h", db_odd.mem_bank[2921],db_even.mem_bank[2921]);
$fdisplay(file, "0x16D40,0x%h_0x%h", db_odd.mem_bank[2922],db_even.mem_bank[2922]);
$fdisplay(file, "0x16D60,0x%h_0x%h", db_odd.mem_bank[2923],db_even.mem_bank[2923]);
$fdisplay(file, "0x16D80,0x%h_0x%h", db_odd.mem_bank[2924],db_even.mem_bank[2924]);
$fdisplay(file, "0x16DA0,0x%h_0x%h", db_odd.mem_bank[2925],db_even.mem_bank[2925]);
$fdisplay(file, "0x16DC0,0x%h_0x%h", db_odd.mem_bank[2926],db_even.mem_bank[2926]);
$fdisplay(file, "0x16DE0,0x%h_0x%h", db_odd.mem_bank[2927],db_even.mem_bank[2927]);
$fdisplay(file, "0x16E00,0x%h_0x%h", db_odd.mem_bank[2928],db_even.mem_bank[2928]);
$fdisplay(file, "0x16E20,0x%h_0x%h", db_odd.mem_bank[2929],db_even.mem_bank[2929]);
$fdisplay(file, "0x16E40,0x%h_0x%h", db_odd.mem_bank[2930],db_even.mem_bank[2930]);
$fdisplay(file, "0x16E60,0x%h_0x%h", db_odd.mem_bank[2931],db_even.mem_bank[2931]);
$fdisplay(file, "0x16E80,0x%h_0x%h", db_odd.mem_bank[2932],db_even.mem_bank[2932]);
$fdisplay(file, "0x16EA0,0x%h_0x%h", db_odd.mem_bank[2933],db_even.mem_bank[2933]);
$fdisplay(file, "0x16EC0,0x%h_0x%h", db_odd.mem_bank[2934],db_even.mem_bank[2934]);
$fdisplay(file, "0x16EE0,0x%h_0x%h", db_odd.mem_bank[2935],db_even.mem_bank[2935]);
$fdisplay(file, "0x16F00,0x%h_0x%h", db_odd.mem_bank[2936],db_even.mem_bank[2936]);
$fdisplay(file, "0x16F20,0x%h_0x%h", db_odd.mem_bank[2937],db_even.mem_bank[2937]);
$fdisplay(file, "0x16F40,0x%h_0x%h", db_odd.mem_bank[2938],db_even.mem_bank[2938]);
$fdisplay(file, "0x16F60,0x%h_0x%h", db_odd.mem_bank[2939],db_even.mem_bank[2939]);
$fdisplay(file, "0x16F80,0x%h_0x%h", db_odd.mem_bank[2940],db_even.mem_bank[2940]);
$fdisplay(file, "0x16FA0,0x%h_0x%h", db_odd.mem_bank[2941],db_even.mem_bank[2941]);
$fdisplay(file, "0x16FC0,0x%h_0x%h", db_odd.mem_bank[2942],db_even.mem_bank[2942]);
$fdisplay(file, "0x16FE0,0x%h_0x%h", db_odd.mem_bank[2943],db_even.mem_bank[2943]);
$fdisplay(file, "0x17000,0x%h_0x%h", db_odd.mem_bank[2944],db_even.mem_bank[2944]);
$fdisplay(file, "0x17020,0x%h_0x%h", db_odd.mem_bank[2945],db_even.mem_bank[2945]);
$fdisplay(file, "0x17040,0x%h_0x%h", db_odd.mem_bank[2946],db_even.mem_bank[2946]);
$fdisplay(file, "0x17060,0x%h_0x%h", db_odd.mem_bank[2947],db_even.mem_bank[2947]);
$fdisplay(file, "0x17080,0x%h_0x%h", db_odd.mem_bank[2948],db_even.mem_bank[2948]);
$fdisplay(file, "0x170A0,0x%h_0x%h", db_odd.mem_bank[2949],db_even.mem_bank[2949]);
$fdisplay(file, "0x170C0,0x%h_0x%h", db_odd.mem_bank[2950],db_even.mem_bank[2950]);
$fdisplay(file, "0x170E0,0x%h_0x%h", db_odd.mem_bank[2951],db_even.mem_bank[2951]);
$fdisplay(file, "0x17100,0x%h_0x%h", db_odd.mem_bank[2952],db_even.mem_bank[2952]);
$fdisplay(file, "0x17120,0x%h_0x%h", db_odd.mem_bank[2953],db_even.mem_bank[2953]);
$fdisplay(file, "0x17140,0x%h_0x%h", db_odd.mem_bank[2954],db_even.mem_bank[2954]);
$fdisplay(file, "0x17160,0x%h_0x%h", db_odd.mem_bank[2955],db_even.mem_bank[2955]);
$fdisplay(file, "0x17180,0x%h_0x%h", db_odd.mem_bank[2956],db_even.mem_bank[2956]);
$fdisplay(file, "0x171A0,0x%h_0x%h", db_odd.mem_bank[2957],db_even.mem_bank[2957]);
$fdisplay(file, "0x171C0,0x%h_0x%h", db_odd.mem_bank[2958],db_even.mem_bank[2958]);
$fdisplay(file, "0x171E0,0x%h_0x%h", db_odd.mem_bank[2959],db_even.mem_bank[2959]);
$fdisplay(file, "0x17200,0x%h_0x%h", db_odd.mem_bank[2960],db_even.mem_bank[2960]);
$fdisplay(file, "0x17220,0x%h_0x%h", db_odd.mem_bank[2961],db_even.mem_bank[2961]);
$fdisplay(file, "0x17240,0x%h_0x%h", db_odd.mem_bank[2962],db_even.mem_bank[2962]);
$fdisplay(file, "0x17260,0x%h_0x%h", db_odd.mem_bank[2963],db_even.mem_bank[2963]);
$fdisplay(file, "0x17280,0x%h_0x%h", db_odd.mem_bank[2964],db_even.mem_bank[2964]);
$fdisplay(file, "0x172A0,0x%h_0x%h", db_odd.mem_bank[2965],db_even.mem_bank[2965]);
$fdisplay(file, "0x172C0,0x%h_0x%h", db_odd.mem_bank[2966],db_even.mem_bank[2966]);
$fdisplay(file, "0x172E0,0x%h_0x%h", db_odd.mem_bank[2967],db_even.mem_bank[2967]);
$fdisplay(file, "0x17300,0x%h_0x%h", db_odd.mem_bank[2968],db_even.mem_bank[2968]);
$fdisplay(file, "0x17320,0x%h_0x%h", db_odd.mem_bank[2969],db_even.mem_bank[2969]);
$fdisplay(file, "0x17340,0x%h_0x%h", db_odd.mem_bank[2970],db_even.mem_bank[2970]);
$fdisplay(file, "0x17360,0x%h_0x%h", db_odd.mem_bank[2971],db_even.mem_bank[2971]);
$fdisplay(file, "0x17380,0x%h_0x%h", db_odd.mem_bank[2972],db_even.mem_bank[2972]);
$fdisplay(file, "0x173A0,0x%h_0x%h", db_odd.mem_bank[2973],db_even.mem_bank[2973]);
$fdisplay(file, "0x173C0,0x%h_0x%h", db_odd.mem_bank[2974],db_even.mem_bank[2974]);
$fdisplay(file, "0x173E0,0x%h_0x%h", db_odd.mem_bank[2975],db_even.mem_bank[2975]);
$fdisplay(file, "0x17400,0x%h_0x%h", db_odd.mem_bank[2976],db_even.mem_bank[2976]);
$fdisplay(file, "0x17420,0x%h_0x%h", db_odd.mem_bank[2977],db_even.mem_bank[2977]);
$fdisplay(file, "0x17440,0x%h_0x%h", db_odd.mem_bank[2978],db_even.mem_bank[2978]);
$fdisplay(file, "0x17460,0x%h_0x%h", db_odd.mem_bank[2979],db_even.mem_bank[2979]);
$fdisplay(file, "0x17480,0x%h_0x%h", db_odd.mem_bank[2980],db_even.mem_bank[2980]);
$fdisplay(file, "0x174A0,0x%h_0x%h", db_odd.mem_bank[2981],db_even.mem_bank[2981]);
$fdisplay(file, "0x174C0,0x%h_0x%h", db_odd.mem_bank[2982],db_even.mem_bank[2982]);
$fdisplay(file, "0x174E0,0x%h_0x%h", db_odd.mem_bank[2983],db_even.mem_bank[2983]);
$fdisplay(file, "0x17500,0x%h_0x%h", db_odd.mem_bank[2984],db_even.mem_bank[2984]);
$fdisplay(file, "0x17520,0x%h_0x%h", db_odd.mem_bank[2985],db_even.mem_bank[2985]);
$fdisplay(file, "0x17540,0x%h_0x%h", db_odd.mem_bank[2986],db_even.mem_bank[2986]);
$fdisplay(file, "0x17560,0x%h_0x%h", db_odd.mem_bank[2987],db_even.mem_bank[2987]);
$fdisplay(file, "0x17580,0x%h_0x%h", db_odd.mem_bank[2988],db_even.mem_bank[2988]);
$fdisplay(file, "0x175A0,0x%h_0x%h", db_odd.mem_bank[2989],db_even.mem_bank[2989]);
$fdisplay(file, "0x175C0,0x%h_0x%h", db_odd.mem_bank[2990],db_even.mem_bank[2990]);
$fdisplay(file, "0x175E0,0x%h_0x%h", db_odd.mem_bank[2991],db_even.mem_bank[2991]);
$fdisplay(file, "0x17600,0x%h_0x%h", db_odd.mem_bank[2992],db_even.mem_bank[2992]);
$fdisplay(file, "0x17620,0x%h_0x%h", db_odd.mem_bank[2993],db_even.mem_bank[2993]);
$fdisplay(file, "0x17640,0x%h_0x%h", db_odd.mem_bank[2994],db_even.mem_bank[2994]);
$fdisplay(file, "0x17660,0x%h_0x%h", db_odd.mem_bank[2995],db_even.mem_bank[2995]);
$fdisplay(file, "0x17680,0x%h_0x%h", db_odd.mem_bank[2996],db_even.mem_bank[2996]);
$fdisplay(file, "0x176A0,0x%h_0x%h", db_odd.mem_bank[2997],db_even.mem_bank[2997]);
$fdisplay(file, "0x176C0,0x%h_0x%h", db_odd.mem_bank[2998],db_even.mem_bank[2998]);
$fdisplay(file, "0x176E0,0x%h_0x%h", db_odd.mem_bank[2999],db_even.mem_bank[2999]);
$fdisplay(file, "0x17700,0x%h_0x%h", db_odd.mem_bank[3000],db_even.mem_bank[3000]);
$fdisplay(file, "0x17720,0x%h_0x%h", db_odd.mem_bank[3001],db_even.mem_bank[3001]);
$fdisplay(file, "0x17740,0x%h_0x%h", db_odd.mem_bank[3002],db_even.mem_bank[3002]);
$fdisplay(file, "0x17760,0x%h_0x%h", db_odd.mem_bank[3003],db_even.mem_bank[3003]);
$fdisplay(file, "0x17780,0x%h_0x%h", db_odd.mem_bank[3004],db_even.mem_bank[3004]);
$fdisplay(file, "0x177A0,0x%h_0x%h", db_odd.mem_bank[3005],db_even.mem_bank[3005]);
$fdisplay(file, "0x177C0,0x%h_0x%h", db_odd.mem_bank[3006],db_even.mem_bank[3006]);
$fdisplay(file, "0x177E0,0x%h_0x%h", db_odd.mem_bank[3007],db_even.mem_bank[3007]);
$fdisplay(file, "0x17800,0x%h_0x%h", db_odd.mem_bank[3008],db_even.mem_bank[3008]);
$fdisplay(file, "0x17820,0x%h_0x%h", db_odd.mem_bank[3009],db_even.mem_bank[3009]);
$fdisplay(file, "0x17840,0x%h_0x%h", db_odd.mem_bank[3010],db_even.mem_bank[3010]);
$fdisplay(file, "0x17860,0x%h_0x%h", db_odd.mem_bank[3011],db_even.mem_bank[3011]);
$fdisplay(file, "0x17880,0x%h_0x%h", db_odd.mem_bank[3012],db_even.mem_bank[3012]);
$fdisplay(file, "0x178A0,0x%h_0x%h", db_odd.mem_bank[3013],db_even.mem_bank[3013]);
$fdisplay(file, "0x178C0,0x%h_0x%h", db_odd.mem_bank[3014],db_even.mem_bank[3014]);
$fdisplay(file, "0x178E0,0x%h_0x%h", db_odd.mem_bank[3015],db_even.mem_bank[3015]);
$fdisplay(file, "0x17900,0x%h_0x%h", db_odd.mem_bank[3016],db_even.mem_bank[3016]);
$fdisplay(file, "0x17920,0x%h_0x%h", db_odd.mem_bank[3017],db_even.mem_bank[3017]);
$fdisplay(file, "0x17940,0x%h_0x%h", db_odd.mem_bank[3018],db_even.mem_bank[3018]);
$fdisplay(file, "0x17960,0x%h_0x%h", db_odd.mem_bank[3019],db_even.mem_bank[3019]);
$fdisplay(file, "0x17980,0x%h_0x%h", db_odd.mem_bank[3020],db_even.mem_bank[3020]);
$fdisplay(file, "0x179A0,0x%h_0x%h", db_odd.mem_bank[3021],db_even.mem_bank[3021]);
$fdisplay(file, "0x179C0,0x%h_0x%h", db_odd.mem_bank[3022],db_even.mem_bank[3022]);
$fdisplay(file, "0x179E0,0x%h_0x%h", db_odd.mem_bank[3023],db_even.mem_bank[3023]);
$fdisplay(file, "0x17A00,0x%h_0x%h", db_odd.mem_bank[3024],db_even.mem_bank[3024]);
$fdisplay(file, "0x17A20,0x%h_0x%h", db_odd.mem_bank[3025],db_even.mem_bank[3025]);
$fdisplay(file, "0x17A40,0x%h_0x%h", db_odd.mem_bank[3026],db_even.mem_bank[3026]);
$fdisplay(file, "0x17A60,0x%h_0x%h", db_odd.mem_bank[3027],db_even.mem_bank[3027]);
$fdisplay(file, "0x17A80,0x%h_0x%h", db_odd.mem_bank[3028],db_even.mem_bank[3028]);
$fdisplay(file, "0x17AA0,0x%h_0x%h", db_odd.mem_bank[3029],db_even.mem_bank[3029]);
$fdisplay(file, "0x17AC0,0x%h_0x%h", db_odd.mem_bank[3030],db_even.mem_bank[3030]);
$fdisplay(file, "0x17AE0,0x%h_0x%h", db_odd.mem_bank[3031],db_even.mem_bank[3031]);
$fdisplay(file, "0x17B00,0x%h_0x%h", db_odd.mem_bank[3032],db_even.mem_bank[3032]);
$fdisplay(file, "0x17B20,0x%h_0x%h", db_odd.mem_bank[3033],db_even.mem_bank[3033]);
$fdisplay(file, "0x17B40,0x%h_0x%h", db_odd.mem_bank[3034],db_even.mem_bank[3034]);
$fdisplay(file, "0x17B60,0x%h_0x%h", db_odd.mem_bank[3035],db_even.mem_bank[3035]);
$fdisplay(file, "0x17B80,0x%h_0x%h", db_odd.mem_bank[3036],db_even.mem_bank[3036]);
$fdisplay(file, "0x17BA0,0x%h_0x%h", db_odd.mem_bank[3037],db_even.mem_bank[3037]);
$fdisplay(file, "0x17BC0,0x%h_0x%h", db_odd.mem_bank[3038],db_even.mem_bank[3038]);
$fdisplay(file, "0x17BE0,0x%h_0x%h", db_odd.mem_bank[3039],db_even.mem_bank[3039]);
$fdisplay(file, "0x17C00,0x%h_0x%h", db_odd.mem_bank[3040],db_even.mem_bank[3040]);
$fdisplay(file, "0x17C20,0x%h_0x%h", db_odd.mem_bank[3041],db_even.mem_bank[3041]);
$fdisplay(file, "0x17C40,0x%h_0x%h", db_odd.mem_bank[3042],db_even.mem_bank[3042]);
$fdisplay(file, "0x17C60,0x%h_0x%h", db_odd.mem_bank[3043],db_even.mem_bank[3043]);
$fdisplay(file, "0x17C80,0x%h_0x%h", db_odd.mem_bank[3044],db_even.mem_bank[3044]);
$fdisplay(file, "0x17CA0,0x%h_0x%h", db_odd.mem_bank[3045],db_even.mem_bank[3045]);
$fdisplay(file, "0x17CC0,0x%h_0x%h", db_odd.mem_bank[3046],db_even.mem_bank[3046]);
$fdisplay(file, "0x17CE0,0x%h_0x%h", db_odd.mem_bank[3047],db_even.mem_bank[3047]);
$fdisplay(file, "0x17D00,0x%h_0x%h", db_odd.mem_bank[3048],db_even.mem_bank[3048]);
$fdisplay(file, "0x17D20,0x%h_0x%h", db_odd.mem_bank[3049],db_even.mem_bank[3049]);
$fdisplay(file, "0x17D40,0x%h_0x%h", db_odd.mem_bank[3050],db_even.mem_bank[3050]);
$fdisplay(file, "0x17D60,0x%h_0x%h", db_odd.mem_bank[3051],db_even.mem_bank[3051]);
$fdisplay(file, "0x17D80,0x%h_0x%h", db_odd.mem_bank[3052],db_even.mem_bank[3052]);
$fdisplay(file, "0x17DA0,0x%h_0x%h", db_odd.mem_bank[3053],db_even.mem_bank[3053]);
$fdisplay(file, "0x17DC0,0x%h_0x%h", db_odd.mem_bank[3054],db_even.mem_bank[3054]);
$fdisplay(file, "0x17DE0,0x%h_0x%h", db_odd.mem_bank[3055],db_even.mem_bank[3055]);
$fdisplay(file, "0x17E00,0x%h_0x%h", db_odd.mem_bank[3056],db_even.mem_bank[3056]);
$fdisplay(file, "0x17E20,0x%h_0x%h", db_odd.mem_bank[3057],db_even.mem_bank[3057]);
$fdisplay(file, "0x17E40,0x%h_0x%h", db_odd.mem_bank[3058],db_even.mem_bank[3058]);
$fdisplay(file, "0x17E60,0x%h_0x%h", db_odd.mem_bank[3059],db_even.mem_bank[3059]);
$fdisplay(file, "0x17E80,0x%h_0x%h", db_odd.mem_bank[3060],db_even.mem_bank[3060]);
$fdisplay(file, "0x17EA0,0x%h_0x%h", db_odd.mem_bank[3061],db_even.mem_bank[3061]);
$fdisplay(file, "0x17EC0,0x%h_0x%h", db_odd.mem_bank[3062],db_even.mem_bank[3062]);
$fdisplay(file, "0x17EE0,0x%h_0x%h", db_odd.mem_bank[3063],db_even.mem_bank[3063]);
$fdisplay(file, "0x17F00,0x%h_0x%h", db_odd.mem_bank[3064],db_even.mem_bank[3064]);
$fdisplay(file, "0x17F20,0x%h_0x%h", db_odd.mem_bank[3065],db_even.mem_bank[3065]);
$fdisplay(file, "0x17F40,0x%h_0x%h", db_odd.mem_bank[3066],db_even.mem_bank[3066]);
$fdisplay(file, "0x17F60,0x%h_0x%h", db_odd.mem_bank[3067],db_even.mem_bank[3067]);
$fdisplay(file, "0x17F80,0x%h_0x%h", db_odd.mem_bank[3068],db_even.mem_bank[3068]);
$fdisplay(file, "0x17FA0,0x%h_0x%h", db_odd.mem_bank[3069],db_even.mem_bank[3069]);
$fdisplay(file, "0x17FC0,0x%h_0x%h", db_odd.mem_bank[3070],db_even.mem_bank[3070]);
$fdisplay(file, "0x17FE0,0x%h_0x%h", db_odd.mem_bank[3071],db_even.mem_bank[3071]);
$fdisplay(file, "0x18000,0x%h_0x%h", db_odd.mem_bank[3072],db_even.mem_bank[3072]);
$fdisplay(file, "0x18020,0x%h_0x%h", db_odd.mem_bank[3073],db_even.mem_bank[3073]);
$fdisplay(file, "0x18040,0x%h_0x%h", db_odd.mem_bank[3074],db_even.mem_bank[3074]);
$fdisplay(file, "0x18060,0x%h_0x%h", db_odd.mem_bank[3075],db_even.mem_bank[3075]);
$fdisplay(file, "0x18080,0x%h_0x%h", db_odd.mem_bank[3076],db_even.mem_bank[3076]);
$fdisplay(file, "0x180A0,0x%h_0x%h", db_odd.mem_bank[3077],db_even.mem_bank[3077]);
$fdisplay(file, "0x180C0,0x%h_0x%h", db_odd.mem_bank[3078],db_even.mem_bank[3078]);
$fdisplay(file, "0x180E0,0x%h_0x%h", db_odd.mem_bank[3079],db_even.mem_bank[3079]);
$fdisplay(file, "0x18100,0x%h_0x%h", db_odd.mem_bank[3080],db_even.mem_bank[3080]);
$fdisplay(file, "0x18120,0x%h_0x%h", db_odd.mem_bank[3081],db_even.mem_bank[3081]);
$fdisplay(file, "0x18140,0x%h_0x%h", db_odd.mem_bank[3082],db_even.mem_bank[3082]);
$fdisplay(file, "0x18160,0x%h_0x%h", db_odd.mem_bank[3083],db_even.mem_bank[3083]);
$fdisplay(file, "0x18180,0x%h_0x%h", db_odd.mem_bank[3084],db_even.mem_bank[3084]);
$fdisplay(file, "0x181A0,0x%h_0x%h", db_odd.mem_bank[3085],db_even.mem_bank[3085]);
$fdisplay(file, "0x181C0,0x%h_0x%h", db_odd.mem_bank[3086],db_even.mem_bank[3086]);
$fdisplay(file, "0x181E0,0x%h_0x%h", db_odd.mem_bank[3087],db_even.mem_bank[3087]);
$fdisplay(file, "0x18200,0x%h_0x%h", db_odd.mem_bank[3088],db_even.mem_bank[3088]);
$fdisplay(file, "0x18220,0x%h_0x%h", db_odd.mem_bank[3089],db_even.mem_bank[3089]);
$fdisplay(file, "0x18240,0x%h_0x%h", db_odd.mem_bank[3090],db_even.mem_bank[3090]);
$fdisplay(file, "0x18260,0x%h_0x%h", db_odd.mem_bank[3091],db_even.mem_bank[3091]);
$fdisplay(file, "0x18280,0x%h_0x%h", db_odd.mem_bank[3092],db_even.mem_bank[3092]);
$fdisplay(file, "0x182A0,0x%h_0x%h", db_odd.mem_bank[3093],db_even.mem_bank[3093]);
$fdisplay(file, "0x182C0,0x%h_0x%h", db_odd.mem_bank[3094],db_even.mem_bank[3094]);
$fdisplay(file, "0x182E0,0x%h_0x%h", db_odd.mem_bank[3095],db_even.mem_bank[3095]);
$fdisplay(file, "0x18300,0x%h_0x%h", db_odd.mem_bank[3096],db_even.mem_bank[3096]);
$fdisplay(file, "0x18320,0x%h_0x%h", db_odd.mem_bank[3097],db_even.mem_bank[3097]);
$fdisplay(file, "0x18340,0x%h_0x%h", db_odd.mem_bank[3098],db_even.mem_bank[3098]);
$fdisplay(file, "0x18360,0x%h_0x%h", db_odd.mem_bank[3099],db_even.mem_bank[3099]);
$fdisplay(file, "0x18380,0x%h_0x%h", db_odd.mem_bank[3100],db_even.mem_bank[3100]);
$fdisplay(file, "0x183A0,0x%h_0x%h", db_odd.mem_bank[3101],db_even.mem_bank[3101]);
$fdisplay(file, "0x183C0,0x%h_0x%h", db_odd.mem_bank[3102],db_even.mem_bank[3102]);
$fdisplay(file, "0x183E0,0x%h_0x%h", db_odd.mem_bank[3103],db_even.mem_bank[3103]);
$fdisplay(file, "0x18400,0x%h_0x%h", db_odd.mem_bank[3104],db_even.mem_bank[3104]);
$fdisplay(file, "0x18420,0x%h_0x%h", db_odd.mem_bank[3105],db_even.mem_bank[3105]);
$fdisplay(file, "0x18440,0x%h_0x%h", db_odd.mem_bank[3106],db_even.mem_bank[3106]);
$fdisplay(file, "0x18460,0x%h_0x%h", db_odd.mem_bank[3107],db_even.mem_bank[3107]);
$fdisplay(file, "0x18480,0x%h_0x%h", db_odd.mem_bank[3108],db_even.mem_bank[3108]);
$fdisplay(file, "0x184A0,0x%h_0x%h", db_odd.mem_bank[3109],db_even.mem_bank[3109]);
$fdisplay(file, "0x184C0,0x%h_0x%h", db_odd.mem_bank[3110],db_even.mem_bank[3110]);
$fdisplay(file, "0x184E0,0x%h_0x%h", db_odd.mem_bank[3111],db_even.mem_bank[3111]);
$fdisplay(file, "0x18500,0x%h_0x%h", db_odd.mem_bank[3112],db_even.mem_bank[3112]);
$fdisplay(file, "0x18520,0x%h_0x%h", db_odd.mem_bank[3113],db_even.mem_bank[3113]);
$fdisplay(file, "0x18540,0x%h_0x%h", db_odd.mem_bank[3114],db_even.mem_bank[3114]);
$fdisplay(file, "0x18560,0x%h_0x%h", db_odd.mem_bank[3115],db_even.mem_bank[3115]);
$fdisplay(file, "0x18580,0x%h_0x%h", db_odd.mem_bank[3116],db_even.mem_bank[3116]);
$fdisplay(file, "0x185A0,0x%h_0x%h", db_odd.mem_bank[3117],db_even.mem_bank[3117]);
$fdisplay(file, "0x185C0,0x%h_0x%h", db_odd.mem_bank[3118],db_even.mem_bank[3118]);
$fdisplay(file, "0x185E0,0x%h_0x%h", db_odd.mem_bank[3119],db_even.mem_bank[3119]);
$fdisplay(file, "0x18600,0x%h_0x%h", db_odd.mem_bank[3120],db_even.mem_bank[3120]);
$fdisplay(file, "0x18620,0x%h_0x%h", db_odd.mem_bank[3121],db_even.mem_bank[3121]);
$fdisplay(file, "0x18640,0x%h_0x%h", db_odd.mem_bank[3122],db_even.mem_bank[3122]);
$fdisplay(file, "0x18660,0x%h_0x%h", db_odd.mem_bank[3123],db_even.mem_bank[3123]);
$fdisplay(file, "0x18680,0x%h_0x%h", db_odd.mem_bank[3124],db_even.mem_bank[3124]);
$fdisplay(file, "0x186A0,0x%h_0x%h", db_odd.mem_bank[3125],db_even.mem_bank[3125]);
$fdisplay(file, "0x186C0,0x%h_0x%h", db_odd.mem_bank[3126],db_even.mem_bank[3126]);
$fdisplay(file, "0x186E0,0x%h_0x%h", db_odd.mem_bank[3127],db_even.mem_bank[3127]);
$fdisplay(file, "0x18700,0x%h_0x%h", db_odd.mem_bank[3128],db_even.mem_bank[3128]);
$fdisplay(file, "0x18720,0x%h_0x%h", db_odd.mem_bank[3129],db_even.mem_bank[3129]);
$fdisplay(file, "0x18740,0x%h_0x%h", db_odd.mem_bank[3130],db_even.mem_bank[3130]);
$fdisplay(file, "0x18760,0x%h_0x%h", db_odd.mem_bank[3131],db_even.mem_bank[3131]);
$fdisplay(file, "0x18780,0x%h_0x%h", db_odd.mem_bank[3132],db_even.mem_bank[3132]);
$fdisplay(file, "0x187A0,0x%h_0x%h", db_odd.mem_bank[3133],db_even.mem_bank[3133]);
$fdisplay(file, "0x187C0,0x%h_0x%h", db_odd.mem_bank[3134],db_even.mem_bank[3134]);
$fdisplay(file, "0x187E0,0x%h_0x%h", db_odd.mem_bank[3135],db_even.mem_bank[3135]);
$fdisplay(file, "0x18800,0x%h_0x%h", db_odd.mem_bank[3136],db_even.mem_bank[3136]);
$fdisplay(file, "0x18820,0x%h_0x%h", db_odd.mem_bank[3137],db_even.mem_bank[3137]);
$fdisplay(file, "0x18840,0x%h_0x%h", db_odd.mem_bank[3138],db_even.mem_bank[3138]);
$fdisplay(file, "0x18860,0x%h_0x%h", db_odd.mem_bank[3139],db_even.mem_bank[3139]);
$fdisplay(file, "0x18880,0x%h_0x%h", db_odd.mem_bank[3140],db_even.mem_bank[3140]);
$fdisplay(file, "0x188A0,0x%h_0x%h", db_odd.mem_bank[3141],db_even.mem_bank[3141]);
$fdisplay(file, "0x188C0,0x%h_0x%h", db_odd.mem_bank[3142],db_even.mem_bank[3142]);
$fdisplay(file, "0x188E0,0x%h_0x%h", db_odd.mem_bank[3143],db_even.mem_bank[3143]);
$fdisplay(file, "0x18900,0x%h_0x%h", db_odd.mem_bank[3144],db_even.mem_bank[3144]);
$fdisplay(file, "0x18920,0x%h_0x%h", db_odd.mem_bank[3145],db_even.mem_bank[3145]);
$fdisplay(file, "0x18940,0x%h_0x%h", db_odd.mem_bank[3146],db_even.mem_bank[3146]);
$fdisplay(file, "0x18960,0x%h_0x%h", db_odd.mem_bank[3147],db_even.mem_bank[3147]);
$fdisplay(file, "0x18980,0x%h_0x%h", db_odd.mem_bank[3148],db_even.mem_bank[3148]);
$fdisplay(file, "0x189A0,0x%h_0x%h", db_odd.mem_bank[3149],db_even.mem_bank[3149]);
$fdisplay(file, "0x189C0,0x%h_0x%h", db_odd.mem_bank[3150],db_even.mem_bank[3150]);
$fdisplay(file, "0x189E0,0x%h_0x%h", db_odd.mem_bank[3151],db_even.mem_bank[3151]);
$fdisplay(file, "0x18A00,0x%h_0x%h", db_odd.mem_bank[3152],db_even.mem_bank[3152]);
$fdisplay(file, "0x18A20,0x%h_0x%h", db_odd.mem_bank[3153],db_even.mem_bank[3153]);
$fdisplay(file, "0x18A40,0x%h_0x%h", db_odd.mem_bank[3154],db_even.mem_bank[3154]);
$fdisplay(file, "0x18A60,0x%h_0x%h", db_odd.mem_bank[3155],db_even.mem_bank[3155]);
$fdisplay(file, "0x18A80,0x%h_0x%h", db_odd.mem_bank[3156],db_even.mem_bank[3156]);
$fdisplay(file, "0x18AA0,0x%h_0x%h", db_odd.mem_bank[3157],db_even.mem_bank[3157]);
$fdisplay(file, "0x18AC0,0x%h_0x%h", db_odd.mem_bank[3158],db_even.mem_bank[3158]);
$fdisplay(file, "0x18AE0,0x%h_0x%h", db_odd.mem_bank[3159],db_even.mem_bank[3159]);
$fdisplay(file, "0x18B00,0x%h_0x%h", db_odd.mem_bank[3160],db_even.mem_bank[3160]);
$fdisplay(file, "0x18B20,0x%h_0x%h", db_odd.mem_bank[3161],db_even.mem_bank[3161]);
$fdisplay(file, "0x18B40,0x%h_0x%h", db_odd.mem_bank[3162],db_even.mem_bank[3162]);
$fdisplay(file, "0x18B60,0x%h_0x%h", db_odd.mem_bank[3163],db_even.mem_bank[3163]);
$fdisplay(file, "0x18B80,0x%h_0x%h", db_odd.mem_bank[3164],db_even.mem_bank[3164]);
$fdisplay(file, "0x18BA0,0x%h_0x%h", db_odd.mem_bank[3165],db_even.mem_bank[3165]);
$fdisplay(file, "0x18BC0,0x%h_0x%h", db_odd.mem_bank[3166],db_even.mem_bank[3166]);
$fdisplay(file, "0x18BE0,0x%h_0x%h", db_odd.mem_bank[3167],db_even.mem_bank[3167]);
$fdisplay(file, "0x18C00,0x%h_0x%h", db_odd.mem_bank[3168],db_even.mem_bank[3168]);
$fdisplay(file, "0x18C20,0x%h_0x%h", db_odd.mem_bank[3169],db_even.mem_bank[3169]);
$fdisplay(file, "0x18C40,0x%h_0x%h", db_odd.mem_bank[3170],db_even.mem_bank[3170]);
$fdisplay(file, "0x18C60,0x%h_0x%h", db_odd.mem_bank[3171],db_even.mem_bank[3171]);
$fdisplay(file, "0x18C80,0x%h_0x%h", db_odd.mem_bank[3172],db_even.mem_bank[3172]);
$fdisplay(file, "0x18CA0,0x%h_0x%h", db_odd.mem_bank[3173],db_even.mem_bank[3173]);
$fdisplay(file, "0x18CC0,0x%h_0x%h", db_odd.mem_bank[3174],db_even.mem_bank[3174]);
$fdisplay(file, "0x18CE0,0x%h_0x%h", db_odd.mem_bank[3175],db_even.mem_bank[3175]);
$fdisplay(file, "0x18D00,0x%h_0x%h", db_odd.mem_bank[3176],db_even.mem_bank[3176]);
$fdisplay(file, "0x18D20,0x%h_0x%h", db_odd.mem_bank[3177],db_even.mem_bank[3177]);
$fdisplay(file, "0x18D40,0x%h_0x%h", db_odd.mem_bank[3178],db_even.mem_bank[3178]);
$fdisplay(file, "0x18D60,0x%h_0x%h", db_odd.mem_bank[3179],db_even.mem_bank[3179]);
$fdisplay(file, "0x18D80,0x%h_0x%h", db_odd.mem_bank[3180],db_even.mem_bank[3180]);
$fdisplay(file, "0x18DA0,0x%h_0x%h", db_odd.mem_bank[3181],db_even.mem_bank[3181]);
$fdisplay(file, "0x18DC0,0x%h_0x%h", db_odd.mem_bank[3182],db_even.mem_bank[3182]);
$fdisplay(file, "0x18DE0,0x%h_0x%h", db_odd.mem_bank[3183],db_even.mem_bank[3183]);
$fdisplay(file, "0x18E00,0x%h_0x%h", db_odd.mem_bank[3184],db_even.mem_bank[3184]);
$fdisplay(file, "0x18E20,0x%h_0x%h", db_odd.mem_bank[3185],db_even.mem_bank[3185]);
$fdisplay(file, "0x18E40,0x%h_0x%h", db_odd.mem_bank[3186],db_even.mem_bank[3186]);
$fdisplay(file, "0x18E60,0x%h_0x%h", db_odd.mem_bank[3187],db_even.mem_bank[3187]);
$fdisplay(file, "0x18E80,0x%h_0x%h", db_odd.mem_bank[3188],db_even.mem_bank[3188]);
$fdisplay(file, "0x18EA0,0x%h_0x%h", db_odd.mem_bank[3189],db_even.mem_bank[3189]);
$fdisplay(file, "0x18EC0,0x%h_0x%h", db_odd.mem_bank[3190],db_even.mem_bank[3190]);
$fdisplay(file, "0x18EE0,0x%h_0x%h", db_odd.mem_bank[3191],db_even.mem_bank[3191]);
$fdisplay(file, "0x18F00,0x%h_0x%h", db_odd.mem_bank[3192],db_even.mem_bank[3192]);
$fdisplay(file, "0x18F20,0x%h_0x%h", db_odd.mem_bank[3193],db_even.mem_bank[3193]);
$fdisplay(file, "0x18F40,0x%h_0x%h", db_odd.mem_bank[3194],db_even.mem_bank[3194]);
$fdisplay(file, "0x18F60,0x%h_0x%h", db_odd.mem_bank[3195],db_even.mem_bank[3195]);
$fdisplay(file, "0x18F80,0x%h_0x%h", db_odd.mem_bank[3196],db_even.mem_bank[3196]);
$fdisplay(file, "0x18FA0,0x%h_0x%h", db_odd.mem_bank[3197],db_even.mem_bank[3197]);
$fdisplay(file, "0x18FC0,0x%h_0x%h", db_odd.mem_bank[3198],db_even.mem_bank[3198]);
$fdisplay(file, "0x18FE0,0x%h_0x%h", db_odd.mem_bank[3199],db_even.mem_bank[3199]);
$fdisplay(file, "0x19000,0x%h_0x%h", db_odd.mem_bank[3200],db_even.mem_bank[3200]);
$fdisplay(file, "0x19020,0x%h_0x%h", db_odd.mem_bank[3201],db_even.mem_bank[3201]);
$fdisplay(file, "0x19040,0x%h_0x%h", db_odd.mem_bank[3202],db_even.mem_bank[3202]);
$fdisplay(file, "0x19060,0x%h_0x%h", db_odd.mem_bank[3203],db_even.mem_bank[3203]);
$fdisplay(file, "0x19080,0x%h_0x%h", db_odd.mem_bank[3204],db_even.mem_bank[3204]);
$fdisplay(file, "0x190A0,0x%h_0x%h", db_odd.mem_bank[3205],db_even.mem_bank[3205]);
$fdisplay(file, "0x190C0,0x%h_0x%h", db_odd.mem_bank[3206],db_even.mem_bank[3206]);
$fdisplay(file, "0x190E0,0x%h_0x%h", db_odd.mem_bank[3207],db_even.mem_bank[3207]);
$fdisplay(file, "0x19100,0x%h_0x%h", db_odd.mem_bank[3208],db_even.mem_bank[3208]);
$fdisplay(file, "0x19120,0x%h_0x%h", db_odd.mem_bank[3209],db_even.mem_bank[3209]);
$fdisplay(file, "0x19140,0x%h_0x%h", db_odd.mem_bank[3210],db_even.mem_bank[3210]);
$fdisplay(file, "0x19160,0x%h_0x%h", db_odd.mem_bank[3211],db_even.mem_bank[3211]);
$fdisplay(file, "0x19180,0x%h_0x%h", db_odd.mem_bank[3212],db_even.mem_bank[3212]);
$fdisplay(file, "0x191A0,0x%h_0x%h", db_odd.mem_bank[3213],db_even.mem_bank[3213]);
$fdisplay(file, "0x191C0,0x%h_0x%h", db_odd.mem_bank[3214],db_even.mem_bank[3214]);
$fdisplay(file, "0x191E0,0x%h_0x%h", db_odd.mem_bank[3215],db_even.mem_bank[3215]);
$fdisplay(file, "0x19200,0x%h_0x%h", db_odd.mem_bank[3216],db_even.mem_bank[3216]);
$fdisplay(file, "0x19220,0x%h_0x%h", db_odd.mem_bank[3217],db_even.mem_bank[3217]);
$fdisplay(file, "0x19240,0x%h_0x%h", db_odd.mem_bank[3218],db_even.mem_bank[3218]);
$fdisplay(file, "0x19260,0x%h_0x%h", db_odd.mem_bank[3219],db_even.mem_bank[3219]);
$fdisplay(file, "0x19280,0x%h_0x%h", db_odd.mem_bank[3220],db_even.mem_bank[3220]);
$fdisplay(file, "0x192A0,0x%h_0x%h", db_odd.mem_bank[3221],db_even.mem_bank[3221]);
$fdisplay(file, "0x192C0,0x%h_0x%h", db_odd.mem_bank[3222],db_even.mem_bank[3222]);
$fdisplay(file, "0x192E0,0x%h_0x%h", db_odd.mem_bank[3223],db_even.mem_bank[3223]);
$fdisplay(file, "0x19300,0x%h_0x%h", db_odd.mem_bank[3224],db_even.mem_bank[3224]);
$fdisplay(file, "0x19320,0x%h_0x%h", db_odd.mem_bank[3225],db_even.mem_bank[3225]);
$fdisplay(file, "0x19340,0x%h_0x%h", db_odd.mem_bank[3226],db_even.mem_bank[3226]);
$fdisplay(file, "0x19360,0x%h_0x%h", db_odd.mem_bank[3227],db_even.mem_bank[3227]);
$fdisplay(file, "0x19380,0x%h_0x%h", db_odd.mem_bank[3228],db_even.mem_bank[3228]);
$fdisplay(file, "0x193A0,0x%h_0x%h", db_odd.mem_bank[3229],db_even.mem_bank[3229]);
$fdisplay(file, "0x193C0,0x%h_0x%h", db_odd.mem_bank[3230],db_even.mem_bank[3230]);
$fdisplay(file, "0x193E0,0x%h_0x%h", db_odd.mem_bank[3231],db_even.mem_bank[3231]);
$fdisplay(file, "0x19400,0x%h_0x%h", db_odd.mem_bank[3232],db_even.mem_bank[3232]);
$fdisplay(file, "0x19420,0x%h_0x%h", db_odd.mem_bank[3233],db_even.mem_bank[3233]);
$fdisplay(file, "0x19440,0x%h_0x%h", db_odd.mem_bank[3234],db_even.mem_bank[3234]);
$fdisplay(file, "0x19460,0x%h_0x%h", db_odd.mem_bank[3235],db_even.mem_bank[3235]);
$fdisplay(file, "0x19480,0x%h_0x%h", db_odd.mem_bank[3236],db_even.mem_bank[3236]);
$fdisplay(file, "0x194A0,0x%h_0x%h", db_odd.mem_bank[3237],db_even.mem_bank[3237]);
$fdisplay(file, "0x194C0,0x%h_0x%h", db_odd.mem_bank[3238],db_even.mem_bank[3238]);
$fdisplay(file, "0x194E0,0x%h_0x%h", db_odd.mem_bank[3239],db_even.mem_bank[3239]);
$fdisplay(file, "0x19500,0x%h_0x%h", db_odd.mem_bank[3240],db_even.mem_bank[3240]);
$fdisplay(file, "0x19520,0x%h_0x%h", db_odd.mem_bank[3241],db_even.mem_bank[3241]);
$fdisplay(file, "0x19540,0x%h_0x%h", db_odd.mem_bank[3242],db_even.mem_bank[3242]);
$fdisplay(file, "0x19560,0x%h_0x%h", db_odd.mem_bank[3243],db_even.mem_bank[3243]);
$fdisplay(file, "0x19580,0x%h_0x%h", db_odd.mem_bank[3244],db_even.mem_bank[3244]);
$fdisplay(file, "0x195A0,0x%h_0x%h", db_odd.mem_bank[3245],db_even.mem_bank[3245]);
$fdisplay(file, "0x195C0,0x%h_0x%h", db_odd.mem_bank[3246],db_even.mem_bank[3246]);
$fdisplay(file, "0x195E0,0x%h_0x%h", db_odd.mem_bank[3247],db_even.mem_bank[3247]);
$fdisplay(file, "0x19600,0x%h_0x%h", db_odd.mem_bank[3248],db_even.mem_bank[3248]);
$fdisplay(file, "0x19620,0x%h_0x%h", db_odd.mem_bank[3249],db_even.mem_bank[3249]);
$fdisplay(file, "0x19640,0x%h_0x%h", db_odd.mem_bank[3250],db_even.mem_bank[3250]);
$fdisplay(file, "0x19660,0x%h_0x%h", db_odd.mem_bank[3251],db_even.mem_bank[3251]);
$fdisplay(file, "0x19680,0x%h_0x%h", db_odd.mem_bank[3252],db_even.mem_bank[3252]);
$fdisplay(file, "0x196A0,0x%h_0x%h", db_odd.mem_bank[3253],db_even.mem_bank[3253]);
$fdisplay(file, "0x196C0,0x%h_0x%h", db_odd.mem_bank[3254],db_even.mem_bank[3254]);
$fdisplay(file, "0x196E0,0x%h_0x%h", db_odd.mem_bank[3255],db_even.mem_bank[3255]);
$fdisplay(file, "0x19700,0x%h_0x%h", db_odd.mem_bank[3256],db_even.mem_bank[3256]);
$fdisplay(file, "0x19720,0x%h_0x%h", db_odd.mem_bank[3257],db_even.mem_bank[3257]);
$fdisplay(file, "0x19740,0x%h_0x%h", db_odd.mem_bank[3258],db_even.mem_bank[3258]);
$fdisplay(file, "0x19760,0x%h_0x%h", db_odd.mem_bank[3259],db_even.mem_bank[3259]);
$fdisplay(file, "0x19780,0x%h_0x%h", db_odd.mem_bank[3260],db_even.mem_bank[3260]);
$fdisplay(file, "0x197A0,0x%h_0x%h", db_odd.mem_bank[3261],db_even.mem_bank[3261]);
$fdisplay(file, "0x197C0,0x%h_0x%h", db_odd.mem_bank[3262],db_even.mem_bank[3262]);
$fdisplay(file, "0x197E0,0x%h_0x%h", db_odd.mem_bank[3263],db_even.mem_bank[3263]);
$fdisplay(file, "0x19800,0x%h_0x%h", db_odd.mem_bank[3264],db_even.mem_bank[3264]);
$fdisplay(file, "0x19820,0x%h_0x%h", db_odd.mem_bank[3265],db_even.mem_bank[3265]);
$fdisplay(file, "0x19840,0x%h_0x%h", db_odd.mem_bank[3266],db_even.mem_bank[3266]);
$fdisplay(file, "0x19860,0x%h_0x%h", db_odd.mem_bank[3267],db_even.mem_bank[3267]);
$fdisplay(file, "0x19880,0x%h_0x%h", db_odd.mem_bank[3268],db_even.mem_bank[3268]);
$fdisplay(file, "0x198A0,0x%h_0x%h", db_odd.mem_bank[3269],db_even.mem_bank[3269]);
$fdisplay(file, "0x198C0,0x%h_0x%h", db_odd.mem_bank[3270],db_even.mem_bank[3270]);
$fdisplay(file, "0x198E0,0x%h_0x%h", db_odd.mem_bank[3271],db_even.mem_bank[3271]);
$fdisplay(file, "0x19900,0x%h_0x%h", db_odd.mem_bank[3272],db_even.mem_bank[3272]);
$fdisplay(file, "0x19920,0x%h_0x%h", db_odd.mem_bank[3273],db_even.mem_bank[3273]);
$fdisplay(file, "0x19940,0x%h_0x%h", db_odd.mem_bank[3274],db_even.mem_bank[3274]);
$fdisplay(file, "0x19960,0x%h_0x%h", db_odd.mem_bank[3275],db_even.mem_bank[3275]);
$fdisplay(file, "0x19980,0x%h_0x%h", db_odd.mem_bank[3276],db_even.mem_bank[3276]);
$fdisplay(file, "0x199A0,0x%h_0x%h", db_odd.mem_bank[3277],db_even.mem_bank[3277]);
$fdisplay(file, "0x199C0,0x%h_0x%h", db_odd.mem_bank[3278],db_even.mem_bank[3278]);
$fdisplay(file, "0x199E0,0x%h_0x%h", db_odd.mem_bank[3279],db_even.mem_bank[3279]);
$fdisplay(file, "0x19A00,0x%h_0x%h", db_odd.mem_bank[3280],db_even.mem_bank[3280]);
$fdisplay(file, "0x19A20,0x%h_0x%h", db_odd.mem_bank[3281],db_even.mem_bank[3281]);
$fdisplay(file, "0x19A40,0x%h_0x%h", db_odd.mem_bank[3282],db_even.mem_bank[3282]);
$fdisplay(file, "0x19A60,0x%h_0x%h", db_odd.mem_bank[3283],db_even.mem_bank[3283]);
$fdisplay(file, "0x19A80,0x%h_0x%h", db_odd.mem_bank[3284],db_even.mem_bank[3284]);
$fdisplay(file, "0x19AA0,0x%h_0x%h", db_odd.mem_bank[3285],db_even.mem_bank[3285]);
$fdisplay(file, "0x19AC0,0x%h_0x%h", db_odd.mem_bank[3286],db_even.mem_bank[3286]);
$fdisplay(file, "0x19AE0,0x%h_0x%h", db_odd.mem_bank[3287],db_even.mem_bank[3287]);
$fdisplay(file, "0x19B00,0x%h_0x%h", db_odd.mem_bank[3288],db_even.mem_bank[3288]);
$fdisplay(file, "0x19B20,0x%h_0x%h", db_odd.mem_bank[3289],db_even.mem_bank[3289]);
$fdisplay(file, "0x19B40,0x%h_0x%h", db_odd.mem_bank[3290],db_even.mem_bank[3290]);
$fdisplay(file, "0x19B60,0x%h_0x%h", db_odd.mem_bank[3291],db_even.mem_bank[3291]);
$fdisplay(file, "0x19B80,0x%h_0x%h", db_odd.mem_bank[3292],db_even.mem_bank[3292]);
$fdisplay(file, "0x19BA0,0x%h_0x%h", db_odd.mem_bank[3293],db_even.mem_bank[3293]);
$fdisplay(file, "0x19BC0,0x%h_0x%h", db_odd.mem_bank[3294],db_even.mem_bank[3294]);
$fdisplay(file, "0x19BE0,0x%h_0x%h", db_odd.mem_bank[3295],db_even.mem_bank[3295]);
$fdisplay(file, "0x19C00,0x%h_0x%h", db_odd.mem_bank[3296],db_even.mem_bank[3296]);
$fdisplay(file, "0x19C20,0x%h_0x%h", db_odd.mem_bank[3297],db_even.mem_bank[3297]);
$fdisplay(file, "0x19C40,0x%h_0x%h", db_odd.mem_bank[3298],db_even.mem_bank[3298]);
$fdisplay(file, "0x19C60,0x%h_0x%h", db_odd.mem_bank[3299],db_even.mem_bank[3299]);
$fdisplay(file, "0x19C80,0x%h_0x%h", db_odd.mem_bank[3300],db_even.mem_bank[3300]);
$fdisplay(file, "0x19CA0,0x%h_0x%h", db_odd.mem_bank[3301],db_even.mem_bank[3301]);
$fdisplay(file, "0x19CC0,0x%h_0x%h", db_odd.mem_bank[3302],db_even.mem_bank[3302]);
$fdisplay(file, "0x19CE0,0x%h_0x%h", db_odd.mem_bank[3303],db_even.mem_bank[3303]);
$fdisplay(file, "0x19D00,0x%h_0x%h", db_odd.mem_bank[3304],db_even.mem_bank[3304]);
$fdisplay(file, "0x19D20,0x%h_0x%h", db_odd.mem_bank[3305],db_even.mem_bank[3305]);
$fdisplay(file, "0x19D40,0x%h_0x%h", db_odd.mem_bank[3306],db_even.mem_bank[3306]);
$fdisplay(file, "0x19D60,0x%h_0x%h", db_odd.mem_bank[3307],db_even.mem_bank[3307]);
$fdisplay(file, "0x19D80,0x%h_0x%h", db_odd.mem_bank[3308],db_even.mem_bank[3308]);
$fdisplay(file, "0x19DA0,0x%h_0x%h", db_odd.mem_bank[3309],db_even.mem_bank[3309]);
$fdisplay(file, "0x19DC0,0x%h_0x%h", db_odd.mem_bank[3310],db_even.mem_bank[3310]);
$fdisplay(file, "0x19DE0,0x%h_0x%h", db_odd.mem_bank[3311],db_even.mem_bank[3311]);
$fdisplay(file, "0x19E00,0x%h_0x%h", db_odd.mem_bank[3312],db_even.mem_bank[3312]);
$fdisplay(file, "0x19E20,0x%h_0x%h", db_odd.mem_bank[3313],db_even.mem_bank[3313]);
$fdisplay(file, "0x19E40,0x%h_0x%h", db_odd.mem_bank[3314],db_even.mem_bank[3314]);
$fdisplay(file, "0x19E60,0x%h_0x%h", db_odd.mem_bank[3315],db_even.mem_bank[3315]);
$fdisplay(file, "0x19E80,0x%h_0x%h", db_odd.mem_bank[3316],db_even.mem_bank[3316]);
$fdisplay(file, "0x19EA0,0x%h_0x%h", db_odd.mem_bank[3317],db_even.mem_bank[3317]);
$fdisplay(file, "0x19EC0,0x%h_0x%h", db_odd.mem_bank[3318],db_even.mem_bank[3318]);
$fdisplay(file, "0x19EE0,0x%h_0x%h", db_odd.mem_bank[3319],db_even.mem_bank[3319]);
$fdisplay(file, "0x19F00,0x%h_0x%h", db_odd.mem_bank[3320],db_even.mem_bank[3320]);
$fdisplay(file, "0x19F20,0x%h_0x%h", db_odd.mem_bank[3321],db_even.mem_bank[3321]);
$fdisplay(file, "0x19F40,0x%h_0x%h", db_odd.mem_bank[3322],db_even.mem_bank[3322]);
$fdisplay(file, "0x19F60,0x%h_0x%h", db_odd.mem_bank[3323],db_even.mem_bank[3323]);
$fdisplay(file, "0x19F80,0x%h_0x%h", db_odd.mem_bank[3324],db_even.mem_bank[3324]);
$fdisplay(file, "0x19FA0,0x%h_0x%h", db_odd.mem_bank[3325],db_even.mem_bank[3325]);
$fdisplay(file, "0x19FC0,0x%h_0x%h", db_odd.mem_bank[3326],db_even.mem_bank[3326]);
$fdisplay(file, "0x19FE0,0x%h_0x%h", db_odd.mem_bank[3327],db_even.mem_bank[3327]);
$fdisplay(file, "0x1A000,0x%h_0x%h", db_odd.mem_bank[3328],db_even.mem_bank[3328]);
$fdisplay(file, "0x1A020,0x%h_0x%h", db_odd.mem_bank[3329],db_even.mem_bank[3329]);
$fdisplay(file, "0x1A040,0x%h_0x%h", db_odd.mem_bank[3330],db_even.mem_bank[3330]);
$fdisplay(file, "0x1A060,0x%h_0x%h", db_odd.mem_bank[3331],db_even.mem_bank[3331]);
$fdisplay(file, "0x1A080,0x%h_0x%h", db_odd.mem_bank[3332],db_even.mem_bank[3332]);
$fdisplay(file, "0x1A0A0,0x%h_0x%h", db_odd.mem_bank[3333],db_even.mem_bank[3333]);
$fdisplay(file, "0x1A0C0,0x%h_0x%h", db_odd.mem_bank[3334],db_even.mem_bank[3334]);
$fdisplay(file, "0x1A0E0,0x%h_0x%h", db_odd.mem_bank[3335],db_even.mem_bank[3335]);
$fdisplay(file, "0x1A100,0x%h_0x%h", db_odd.mem_bank[3336],db_even.mem_bank[3336]);
$fdisplay(file, "0x1A120,0x%h_0x%h", db_odd.mem_bank[3337],db_even.mem_bank[3337]);
$fdisplay(file, "0x1A140,0x%h_0x%h", db_odd.mem_bank[3338],db_even.mem_bank[3338]);
$fdisplay(file, "0x1A160,0x%h_0x%h", db_odd.mem_bank[3339],db_even.mem_bank[3339]);
$fdisplay(file, "0x1A180,0x%h_0x%h", db_odd.mem_bank[3340],db_even.mem_bank[3340]);
$fdisplay(file, "0x1A1A0,0x%h_0x%h", db_odd.mem_bank[3341],db_even.mem_bank[3341]);
$fdisplay(file, "0x1A1C0,0x%h_0x%h", db_odd.mem_bank[3342],db_even.mem_bank[3342]);
$fdisplay(file, "0x1A1E0,0x%h_0x%h", db_odd.mem_bank[3343],db_even.mem_bank[3343]);
$fdisplay(file, "0x1A200,0x%h_0x%h", db_odd.mem_bank[3344],db_even.mem_bank[3344]);
$fdisplay(file, "0x1A220,0x%h_0x%h", db_odd.mem_bank[3345],db_even.mem_bank[3345]);
$fdisplay(file, "0x1A240,0x%h_0x%h", db_odd.mem_bank[3346],db_even.mem_bank[3346]);
$fdisplay(file, "0x1A260,0x%h_0x%h", db_odd.mem_bank[3347],db_even.mem_bank[3347]);
$fdisplay(file, "0x1A280,0x%h_0x%h", db_odd.mem_bank[3348],db_even.mem_bank[3348]);
$fdisplay(file, "0x1A2A0,0x%h_0x%h", db_odd.mem_bank[3349],db_even.mem_bank[3349]);
$fdisplay(file, "0x1A2C0,0x%h_0x%h", db_odd.mem_bank[3350],db_even.mem_bank[3350]);
$fdisplay(file, "0x1A2E0,0x%h_0x%h", db_odd.mem_bank[3351],db_even.mem_bank[3351]);
$fdisplay(file, "0x1A300,0x%h_0x%h", db_odd.mem_bank[3352],db_even.mem_bank[3352]);
$fdisplay(file, "0x1A320,0x%h_0x%h", db_odd.mem_bank[3353],db_even.mem_bank[3353]);
$fdisplay(file, "0x1A340,0x%h_0x%h", db_odd.mem_bank[3354],db_even.mem_bank[3354]);
$fdisplay(file, "0x1A360,0x%h_0x%h", db_odd.mem_bank[3355],db_even.mem_bank[3355]);
$fdisplay(file, "0x1A380,0x%h_0x%h", db_odd.mem_bank[3356],db_even.mem_bank[3356]);
$fdisplay(file, "0x1A3A0,0x%h_0x%h", db_odd.mem_bank[3357],db_even.mem_bank[3357]);
$fdisplay(file, "0x1A3C0,0x%h_0x%h", db_odd.mem_bank[3358],db_even.mem_bank[3358]);
$fdisplay(file, "0x1A3E0,0x%h_0x%h", db_odd.mem_bank[3359],db_even.mem_bank[3359]);
$fdisplay(file, "0x1A400,0x%h_0x%h", db_odd.mem_bank[3360],db_even.mem_bank[3360]);
$fdisplay(file, "0x1A420,0x%h_0x%h", db_odd.mem_bank[3361],db_even.mem_bank[3361]);
$fdisplay(file, "0x1A440,0x%h_0x%h", db_odd.mem_bank[3362],db_even.mem_bank[3362]);
$fdisplay(file, "0x1A460,0x%h_0x%h", db_odd.mem_bank[3363],db_even.mem_bank[3363]);
$fdisplay(file, "0x1A480,0x%h_0x%h", db_odd.mem_bank[3364],db_even.mem_bank[3364]);
$fdisplay(file, "0x1A4A0,0x%h_0x%h", db_odd.mem_bank[3365],db_even.mem_bank[3365]);
$fdisplay(file, "0x1A4C0,0x%h_0x%h", db_odd.mem_bank[3366],db_even.mem_bank[3366]);
$fdisplay(file, "0x1A4E0,0x%h_0x%h", db_odd.mem_bank[3367],db_even.mem_bank[3367]);
$fdisplay(file, "0x1A500,0x%h_0x%h", db_odd.mem_bank[3368],db_even.mem_bank[3368]);
$fdisplay(file, "0x1A520,0x%h_0x%h", db_odd.mem_bank[3369],db_even.mem_bank[3369]);
$fdisplay(file, "0x1A540,0x%h_0x%h", db_odd.mem_bank[3370],db_even.mem_bank[3370]);
$fdisplay(file, "0x1A560,0x%h_0x%h", db_odd.mem_bank[3371],db_even.mem_bank[3371]);
$fdisplay(file, "0x1A580,0x%h_0x%h", db_odd.mem_bank[3372],db_even.mem_bank[3372]);
$fdisplay(file, "0x1A5A0,0x%h_0x%h", db_odd.mem_bank[3373],db_even.mem_bank[3373]);
$fdisplay(file, "0x1A5C0,0x%h_0x%h", db_odd.mem_bank[3374],db_even.mem_bank[3374]);
$fdisplay(file, "0x1A5E0,0x%h_0x%h", db_odd.mem_bank[3375],db_even.mem_bank[3375]);
$fdisplay(file, "0x1A600,0x%h_0x%h", db_odd.mem_bank[3376],db_even.mem_bank[3376]);
$fdisplay(file, "0x1A620,0x%h_0x%h", db_odd.mem_bank[3377],db_even.mem_bank[3377]);
$fdisplay(file, "0x1A640,0x%h_0x%h", db_odd.mem_bank[3378],db_even.mem_bank[3378]);
$fdisplay(file, "0x1A660,0x%h_0x%h", db_odd.mem_bank[3379],db_even.mem_bank[3379]);
$fdisplay(file, "0x1A680,0x%h_0x%h", db_odd.mem_bank[3380],db_even.mem_bank[3380]);
$fdisplay(file, "0x1A6A0,0x%h_0x%h", db_odd.mem_bank[3381],db_even.mem_bank[3381]);
$fdisplay(file, "0x1A6C0,0x%h_0x%h", db_odd.mem_bank[3382],db_even.mem_bank[3382]);
$fdisplay(file, "0x1A6E0,0x%h_0x%h", db_odd.mem_bank[3383],db_even.mem_bank[3383]);
$fdisplay(file, "0x1A700,0x%h_0x%h", db_odd.mem_bank[3384],db_even.mem_bank[3384]);
$fdisplay(file, "0x1A720,0x%h_0x%h", db_odd.mem_bank[3385],db_even.mem_bank[3385]);
$fdisplay(file, "0x1A740,0x%h_0x%h", db_odd.mem_bank[3386],db_even.mem_bank[3386]);
$fdisplay(file, "0x1A760,0x%h_0x%h", db_odd.mem_bank[3387],db_even.mem_bank[3387]);
$fdisplay(file, "0x1A780,0x%h_0x%h", db_odd.mem_bank[3388],db_even.mem_bank[3388]);
$fdisplay(file, "0x1A7A0,0x%h_0x%h", db_odd.mem_bank[3389],db_even.mem_bank[3389]);
$fdisplay(file, "0x1A7C0,0x%h_0x%h", db_odd.mem_bank[3390],db_even.mem_bank[3390]);
$fdisplay(file, "0x1A7E0,0x%h_0x%h", db_odd.mem_bank[3391],db_even.mem_bank[3391]);
$fdisplay(file, "0x1A800,0x%h_0x%h", db_odd.mem_bank[3392],db_even.mem_bank[3392]);
$fdisplay(file, "0x1A820,0x%h_0x%h", db_odd.mem_bank[3393],db_even.mem_bank[3393]);
$fdisplay(file, "0x1A840,0x%h_0x%h", db_odd.mem_bank[3394],db_even.mem_bank[3394]);
$fdisplay(file, "0x1A860,0x%h_0x%h", db_odd.mem_bank[3395],db_even.mem_bank[3395]);
$fdisplay(file, "0x1A880,0x%h_0x%h", db_odd.mem_bank[3396],db_even.mem_bank[3396]);
$fdisplay(file, "0x1A8A0,0x%h_0x%h", db_odd.mem_bank[3397],db_even.mem_bank[3397]);
$fdisplay(file, "0x1A8C0,0x%h_0x%h", db_odd.mem_bank[3398],db_even.mem_bank[3398]);
$fdisplay(file, "0x1A8E0,0x%h_0x%h", db_odd.mem_bank[3399],db_even.mem_bank[3399]);
$fdisplay(file, "0x1A900,0x%h_0x%h", db_odd.mem_bank[3400],db_even.mem_bank[3400]);
$fdisplay(file, "0x1A920,0x%h_0x%h", db_odd.mem_bank[3401],db_even.mem_bank[3401]);
$fdisplay(file, "0x1A940,0x%h_0x%h", db_odd.mem_bank[3402],db_even.mem_bank[3402]);
$fdisplay(file, "0x1A960,0x%h_0x%h", db_odd.mem_bank[3403],db_even.mem_bank[3403]);
$fdisplay(file, "0x1A980,0x%h_0x%h", db_odd.mem_bank[3404],db_even.mem_bank[3404]);
$fdisplay(file, "0x1A9A0,0x%h_0x%h", db_odd.mem_bank[3405],db_even.mem_bank[3405]);
$fdisplay(file, "0x1A9C0,0x%h_0x%h", db_odd.mem_bank[3406],db_even.mem_bank[3406]);
$fdisplay(file, "0x1A9E0,0x%h_0x%h", db_odd.mem_bank[3407],db_even.mem_bank[3407]);
$fdisplay(file, "0x1AA00,0x%h_0x%h", db_odd.mem_bank[3408],db_even.mem_bank[3408]);
$fdisplay(file, "0x1AA20,0x%h_0x%h", db_odd.mem_bank[3409],db_even.mem_bank[3409]);
$fdisplay(file, "0x1AA40,0x%h_0x%h", db_odd.mem_bank[3410],db_even.mem_bank[3410]);
$fdisplay(file, "0x1AA60,0x%h_0x%h", db_odd.mem_bank[3411],db_even.mem_bank[3411]);
$fdisplay(file, "0x1AA80,0x%h_0x%h", db_odd.mem_bank[3412],db_even.mem_bank[3412]);
$fdisplay(file, "0x1AAA0,0x%h_0x%h", db_odd.mem_bank[3413],db_even.mem_bank[3413]);
$fdisplay(file, "0x1AAC0,0x%h_0x%h", db_odd.mem_bank[3414],db_even.mem_bank[3414]);
$fdisplay(file, "0x1AAE0,0x%h_0x%h", db_odd.mem_bank[3415],db_even.mem_bank[3415]);
$fdisplay(file, "0x1AB00,0x%h_0x%h", db_odd.mem_bank[3416],db_even.mem_bank[3416]);
$fdisplay(file, "0x1AB20,0x%h_0x%h", db_odd.mem_bank[3417],db_even.mem_bank[3417]);
$fdisplay(file, "0x1AB40,0x%h_0x%h", db_odd.mem_bank[3418],db_even.mem_bank[3418]);
$fdisplay(file, "0x1AB60,0x%h_0x%h", db_odd.mem_bank[3419],db_even.mem_bank[3419]);
$fdisplay(file, "0x1AB80,0x%h_0x%h", db_odd.mem_bank[3420],db_even.mem_bank[3420]);
$fdisplay(file, "0x1ABA0,0x%h_0x%h", db_odd.mem_bank[3421],db_even.mem_bank[3421]);
$fdisplay(file, "0x1ABC0,0x%h_0x%h", db_odd.mem_bank[3422],db_even.mem_bank[3422]);
$fdisplay(file, "0x1ABE0,0x%h_0x%h", db_odd.mem_bank[3423],db_even.mem_bank[3423]);
$fdisplay(file, "0x1AC00,0x%h_0x%h", db_odd.mem_bank[3424],db_even.mem_bank[3424]);
$fdisplay(file, "0x1AC20,0x%h_0x%h", db_odd.mem_bank[3425],db_even.mem_bank[3425]);
$fdisplay(file, "0x1AC40,0x%h_0x%h", db_odd.mem_bank[3426],db_even.mem_bank[3426]);
$fdisplay(file, "0x1AC60,0x%h_0x%h", db_odd.mem_bank[3427],db_even.mem_bank[3427]);
$fdisplay(file, "0x1AC80,0x%h_0x%h", db_odd.mem_bank[3428],db_even.mem_bank[3428]);
$fdisplay(file, "0x1ACA0,0x%h_0x%h", db_odd.mem_bank[3429],db_even.mem_bank[3429]);
$fdisplay(file, "0x1ACC0,0x%h_0x%h", db_odd.mem_bank[3430],db_even.mem_bank[3430]);
$fdisplay(file, "0x1ACE0,0x%h_0x%h", db_odd.mem_bank[3431],db_even.mem_bank[3431]);
$fdisplay(file, "0x1AD00,0x%h_0x%h", db_odd.mem_bank[3432],db_even.mem_bank[3432]);
$fdisplay(file, "0x1AD20,0x%h_0x%h", db_odd.mem_bank[3433],db_even.mem_bank[3433]);
$fdisplay(file, "0x1AD40,0x%h_0x%h", db_odd.mem_bank[3434],db_even.mem_bank[3434]);
$fdisplay(file, "0x1AD60,0x%h_0x%h", db_odd.mem_bank[3435],db_even.mem_bank[3435]);
$fdisplay(file, "0x1AD80,0x%h_0x%h", db_odd.mem_bank[3436],db_even.mem_bank[3436]);
$fdisplay(file, "0x1ADA0,0x%h_0x%h", db_odd.mem_bank[3437],db_even.mem_bank[3437]);
$fdisplay(file, "0x1ADC0,0x%h_0x%h", db_odd.mem_bank[3438],db_even.mem_bank[3438]);
$fdisplay(file, "0x1ADE0,0x%h_0x%h", db_odd.mem_bank[3439],db_even.mem_bank[3439]);
$fdisplay(file, "0x1AE00,0x%h_0x%h", db_odd.mem_bank[3440],db_even.mem_bank[3440]);
$fdisplay(file, "0x1AE20,0x%h_0x%h", db_odd.mem_bank[3441],db_even.mem_bank[3441]);
$fdisplay(file, "0x1AE40,0x%h_0x%h", db_odd.mem_bank[3442],db_even.mem_bank[3442]);
$fdisplay(file, "0x1AE60,0x%h_0x%h", db_odd.mem_bank[3443],db_even.mem_bank[3443]);
$fdisplay(file, "0x1AE80,0x%h_0x%h", db_odd.mem_bank[3444],db_even.mem_bank[3444]);
$fdisplay(file, "0x1AEA0,0x%h_0x%h", db_odd.mem_bank[3445],db_even.mem_bank[3445]);
$fdisplay(file, "0x1AEC0,0x%h_0x%h", db_odd.mem_bank[3446],db_even.mem_bank[3446]);
$fdisplay(file, "0x1AEE0,0x%h_0x%h", db_odd.mem_bank[3447],db_even.mem_bank[3447]);
$fdisplay(file, "0x1AF00,0x%h_0x%h", db_odd.mem_bank[3448],db_even.mem_bank[3448]);
$fdisplay(file, "0x1AF20,0x%h_0x%h", db_odd.mem_bank[3449],db_even.mem_bank[3449]);
$fdisplay(file, "0x1AF40,0x%h_0x%h", db_odd.mem_bank[3450],db_even.mem_bank[3450]);
$fdisplay(file, "0x1AF60,0x%h_0x%h", db_odd.mem_bank[3451],db_even.mem_bank[3451]);
$fdisplay(file, "0x1AF80,0x%h_0x%h", db_odd.mem_bank[3452],db_even.mem_bank[3452]);
$fdisplay(file, "0x1AFA0,0x%h_0x%h", db_odd.mem_bank[3453],db_even.mem_bank[3453]);
$fdisplay(file, "0x1AFC0,0x%h_0x%h", db_odd.mem_bank[3454],db_even.mem_bank[3454]);
$fdisplay(file, "0x1AFE0,0x%h_0x%h", db_odd.mem_bank[3455],db_even.mem_bank[3455]);
$fdisplay(file, "0x1B000,0x%h_0x%h", db_odd.mem_bank[3456],db_even.mem_bank[3456]);
$fdisplay(file, "0x1B020,0x%h_0x%h", db_odd.mem_bank[3457],db_even.mem_bank[3457]);
$fdisplay(file, "0x1B040,0x%h_0x%h", db_odd.mem_bank[3458],db_even.mem_bank[3458]);
$fdisplay(file, "0x1B060,0x%h_0x%h", db_odd.mem_bank[3459],db_even.mem_bank[3459]);
$fdisplay(file, "0x1B080,0x%h_0x%h", db_odd.mem_bank[3460],db_even.mem_bank[3460]);
$fdisplay(file, "0x1B0A0,0x%h_0x%h", db_odd.mem_bank[3461],db_even.mem_bank[3461]);
$fdisplay(file, "0x1B0C0,0x%h_0x%h", db_odd.mem_bank[3462],db_even.mem_bank[3462]);
$fdisplay(file, "0x1B0E0,0x%h_0x%h", db_odd.mem_bank[3463],db_even.mem_bank[3463]);
$fdisplay(file, "0x1B100,0x%h_0x%h", db_odd.mem_bank[3464],db_even.mem_bank[3464]);
$fdisplay(file, "0x1B120,0x%h_0x%h", db_odd.mem_bank[3465],db_even.mem_bank[3465]);
$fdisplay(file, "0x1B140,0x%h_0x%h", db_odd.mem_bank[3466],db_even.mem_bank[3466]);
$fdisplay(file, "0x1B160,0x%h_0x%h", db_odd.mem_bank[3467],db_even.mem_bank[3467]);
$fdisplay(file, "0x1B180,0x%h_0x%h", db_odd.mem_bank[3468],db_even.mem_bank[3468]);
$fdisplay(file, "0x1B1A0,0x%h_0x%h", db_odd.mem_bank[3469],db_even.mem_bank[3469]);
$fdisplay(file, "0x1B1C0,0x%h_0x%h", db_odd.mem_bank[3470],db_even.mem_bank[3470]);
$fdisplay(file, "0x1B1E0,0x%h_0x%h", db_odd.mem_bank[3471],db_even.mem_bank[3471]);
$fdisplay(file, "0x1B200,0x%h_0x%h", db_odd.mem_bank[3472],db_even.mem_bank[3472]);
$fdisplay(file, "0x1B220,0x%h_0x%h", db_odd.mem_bank[3473],db_even.mem_bank[3473]);
$fdisplay(file, "0x1B240,0x%h_0x%h", db_odd.mem_bank[3474],db_even.mem_bank[3474]);
$fdisplay(file, "0x1B260,0x%h_0x%h", db_odd.mem_bank[3475],db_even.mem_bank[3475]);
$fdisplay(file, "0x1B280,0x%h_0x%h", db_odd.mem_bank[3476],db_even.mem_bank[3476]);
$fdisplay(file, "0x1B2A0,0x%h_0x%h", db_odd.mem_bank[3477],db_even.mem_bank[3477]);
$fdisplay(file, "0x1B2C0,0x%h_0x%h", db_odd.mem_bank[3478],db_even.mem_bank[3478]);
$fdisplay(file, "0x1B2E0,0x%h_0x%h", db_odd.mem_bank[3479],db_even.mem_bank[3479]);
$fdisplay(file, "0x1B300,0x%h_0x%h", db_odd.mem_bank[3480],db_even.mem_bank[3480]);
$fdisplay(file, "0x1B320,0x%h_0x%h", db_odd.mem_bank[3481],db_even.mem_bank[3481]);
$fdisplay(file, "0x1B340,0x%h_0x%h", db_odd.mem_bank[3482],db_even.mem_bank[3482]);
$fdisplay(file, "0x1B360,0x%h_0x%h", db_odd.mem_bank[3483],db_even.mem_bank[3483]);
$fdisplay(file, "0x1B380,0x%h_0x%h", db_odd.mem_bank[3484],db_even.mem_bank[3484]);
$fdisplay(file, "0x1B3A0,0x%h_0x%h", db_odd.mem_bank[3485],db_even.mem_bank[3485]);
$fdisplay(file, "0x1B3C0,0x%h_0x%h", db_odd.mem_bank[3486],db_even.mem_bank[3486]);
$fdisplay(file, "0x1B3E0,0x%h_0x%h", db_odd.mem_bank[3487],db_even.mem_bank[3487]);
$fdisplay(file, "0x1B400,0x%h_0x%h", db_odd.mem_bank[3488],db_even.mem_bank[3488]);
$fdisplay(file, "0x1B420,0x%h_0x%h", db_odd.mem_bank[3489],db_even.mem_bank[3489]);
$fdisplay(file, "0x1B440,0x%h_0x%h", db_odd.mem_bank[3490],db_even.mem_bank[3490]);
$fdisplay(file, "0x1B460,0x%h_0x%h", db_odd.mem_bank[3491],db_even.mem_bank[3491]);
$fdisplay(file, "0x1B480,0x%h_0x%h", db_odd.mem_bank[3492],db_even.mem_bank[3492]);
$fdisplay(file, "0x1B4A0,0x%h_0x%h", db_odd.mem_bank[3493],db_even.mem_bank[3493]);
$fdisplay(file, "0x1B4C0,0x%h_0x%h", db_odd.mem_bank[3494],db_even.mem_bank[3494]);
$fdisplay(file, "0x1B4E0,0x%h_0x%h", db_odd.mem_bank[3495],db_even.mem_bank[3495]);
$fdisplay(file, "0x1B500,0x%h_0x%h", db_odd.mem_bank[3496],db_even.mem_bank[3496]);
$fdisplay(file, "0x1B520,0x%h_0x%h", db_odd.mem_bank[3497],db_even.mem_bank[3497]);
$fdisplay(file, "0x1B540,0x%h_0x%h", db_odd.mem_bank[3498],db_even.mem_bank[3498]);
$fdisplay(file, "0x1B560,0x%h_0x%h", db_odd.mem_bank[3499],db_even.mem_bank[3499]);
$fdisplay(file, "0x1B580,0x%h_0x%h", db_odd.mem_bank[3500],db_even.mem_bank[3500]);
$fdisplay(file, "0x1B5A0,0x%h_0x%h", db_odd.mem_bank[3501],db_even.mem_bank[3501]);
$fdisplay(file, "0x1B5C0,0x%h_0x%h", db_odd.mem_bank[3502],db_even.mem_bank[3502]);
$fdisplay(file, "0x1B5E0,0x%h_0x%h", db_odd.mem_bank[3503],db_even.mem_bank[3503]);
$fdisplay(file, "0x1B600,0x%h_0x%h", db_odd.mem_bank[3504],db_even.mem_bank[3504]);
$fdisplay(file, "0x1B620,0x%h_0x%h", db_odd.mem_bank[3505],db_even.mem_bank[3505]);
$fdisplay(file, "0x1B640,0x%h_0x%h", db_odd.mem_bank[3506],db_even.mem_bank[3506]);
$fdisplay(file, "0x1B660,0x%h_0x%h", db_odd.mem_bank[3507],db_even.mem_bank[3507]);
$fdisplay(file, "0x1B680,0x%h_0x%h", db_odd.mem_bank[3508],db_even.mem_bank[3508]);
$fdisplay(file, "0x1B6A0,0x%h_0x%h", db_odd.mem_bank[3509],db_even.mem_bank[3509]);
$fdisplay(file, "0x1B6C0,0x%h_0x%h", db_odd.mem_bank[3510],db_even.mem_bank[3510]);
$fdisplay(file, "0x1B6E0,0x%h_0x%h", db_odd.mem_bank[3511],db_even.mem_bank[3511]);
$fdisplay(file, "0x1B700,0x%h_0x%h", db_odd.mem_bank[3512],db_even.mem_bank[3512]);
$fdisplay(file, "0x1B720,0x%h_0x%h", db_odd.mem_bank[3513],db_even.mem_bank[3513]);
$fdisplay(file, "0x1B740,0x%h_0x%h", db_odd.mem_bank[3514],db_even.mem_bank[3514]);
$fdisplay(file, "0x1B760,0x%h_0x%h", db_odd.mem_bank[3515],db_even.mem_bank[3515]);
$fdisplay(file, "0x1B780,0x%h_0x%h", db_odd.mem_bank[3516],db_even.mem_bank[3516]);
$fdisplay(file, "0x1B7A0,0x%h_0x%h", db_odd.mem_bank[3517],db_even.mem_bank[3517]);
$fdisplay(file, "0x1B7C0,0x%h_0x%h", db_odd.mem_bank[3518],db_even.mem_bank[3518]);
$fdisplay(file, "0x1B7E0,0x%h_0x%h", db_odd.mem_bank[3519],db_even.mem_bank[3519]);
$fdisplay(file, "0x1B800,0x%h_0x%h", db_odd.mem_bank[3520],db_even.mem_bank[3520]);
$fdisplay(file, "0x1B820,0x%h_0x%h", db_odd.mem_bank[3521],db_even.mem_bank[3521]);
$fdisplay(file, "0x1B840,0x%h_0x%h", db_odd.mem_bank[3522],db_even.mem_bank[3522]);
$fdisplay(file, "0x1B860,0x%h_0x%h", db_odd.mem_bank[3523],db_even.mem_bank[3523]);
$fdisplay(file, "0x1B880,0x%h_0x%h", db_odd.mem_bank[3524],db_even.mem_bank[3524]);
$fdisplay(file, "0x1B8A0,0x%h_0x%h", db_odd.mem_bank[3525],db_even.mem_bank[3525]);
$fdisplay(file, "0x1B8C0,0x%h_0x%h", db_odd.mem_bank[3526],db_even.mem_bank[3526]);
$fdisplay(file, "0x1B8E0,0x%h_0x%h", db_odd.mem_bank[3527],db_even.mem_bank[3527]);
$fdisplay(file, "0x1B900,0x%h_0x%h", db_odd.mem_bank[3528],db_even.mem_bank[3528]);
$fdisplay(file, "0x1B920,0x%h_0x%h", db_odd.mem_bank[3529],db_even.mem_bank[3529]);
$fdisplay(file, "0x1B940,0x%h_0x%h", db_odd.mem_bank[3530],db_even.mem_bank[3530]);
$fdisplay(file, "0x1B960,0x%h_0x%h", db_odd.mem_bank[3531],db_even.mem_bank[3531]);
$fdisplay(file, "0x1B980,0x%h_0x%h", db_odd.mem_bank[3532],db_even.mem_bank[3532]);
$fdisplay(file, "0x1B9A0,0x%h_0x%h", db_odd.mem_bank[3533],db_even.mem_bank[3533]);
$fdisplay(file, "0x1B9C0,0x%h_0x%h", db_odd.mem_bank[3534],db_even.mem_bank[3534]);
$fdisplay(file, "0x1B9E0,0x%h_0x%h", db_odd.mem_bank[3535],db_even.mem_bank[3535]);
$fdisplay(file, "0x1BA00,0x%h_0x%h", db_odd.mem_bank[3536],db_even.mem_bank[3536]);
$fdisplay(file, "0x1BA20,0x%h_0x%h", db_odd.mem_bank[3537],db_even.mem_bank[3537]);
$fdisplay(file, "0x1BA40,0x%h_0x%h", db_odd.mem_bank[3538],db_even.mem_bank[3538]);
$fdisplay(file, "0x1BA60,0x%h_0x%h", db_odd.mem_bank[3539],db_even.mem_bank[3539]);
$fdisplay(file, "0x1BA80,0x%h_0x%h", db_odd.mem_bank[3540],db_even.mem_bank[3540]);
$fdisplay(file, "0x1BAA0,0x%h_0x%h", db_odd.mem_bank[3541],db_even.mem_bank[3541]);
$fdisplay(file, "0x1BAC0,0x%h_0x%h", db_odd.mem_bank[3542],db_even.mem_bank[3542]);
$fdisplay(file, "0x1BAE0,0x%h_0x%h", db_odd.mem_bank[3543],db_even.mem_bank[3543]);
$fdisplay(file, "0x1BB00,0x%h_0x%h", db_odd.mem_bank[3544],db_even.mem_bank[3544]);
$fdisplay(file, "0x1BB20,0x%h_0x%h", db_odd.mem_bank[3545],db_even.mem_bank[3545]);
$fdisplay(file, "0x1BB40,0x%h_0x%h", db_odd.mem_bank[3546],db_even.mem_bank[3546]);
$fdisplay(file, "0x1BB60,0x%h_0x%h", db_odd.mem_bank[3547],db_even.mem_bank[3547]);
$fdisplay(file, "0x1BB80,0x%h_0x%h", db_odd.mem_bank[3548],db_even.mem_bank[3548]);
$fdisplay(file, "0x1BBA0,0x%h_0x%h", db_odd.mem_bank[3549],db_even.mem_bank[3549]);
$fdisplay(file, "0x1BBC0,0x%h_0x%h", db_odd.mem_bank[3550],db_even.mem_bank[3550]);
$fdisplay(file, "0x1BBE0,0x%h_0x%h", db_odd.mem_bank[3551],db_even.mem_bank[3551]);
$fdisplay(file, "0x1BC00,0x%h_0x%h", db_odd.mem_bank[3552],db_even.mem_bank[3552]);
$fdisplay(file, "0x1BC20,0x%h_0x%h", db_odd.mem_bank[3553],db_even.mem_bank[3553]);
$fdisplay(file, "0x1BC40,0x%h_0x%h", db_odd.mem_bank[3554],db_even.mem_bank[3554]);
$fdisplay(file, "0x1BC60,0x%h_0x%h", db_odd.mem_bank[3555],db_even.mem_bank[3555]);
$fdisplay(file, "0x1BC80,0x%h_0x%h", db_odd.mem_bank[3556],db_even.mem_bank[3556]);
$fdisplay(file, "0x1BCA0,0x%h_0x%h", db_odd.mem_bank[3557],db_even.mem_bank[3557]);
$fdisplay(file, "0x1BCC0,0x%h_0x%h", db_odd.mem_bank[3558],db_even.mem_bank[3558]);
$fdisplay(file, "0x1BCE0,0x%h_0x%h", db_odd.mem_bank[3559],db_even.mem_bank[3559]);
$fdisplay(file, "0x1BD00,0x%h_0x%h", db_odd.mem_bank[3560],db_even.mem_bank[3560]);
$fdisplay(file, "0x1BD20,0x%h_0x%h", db_odd.mem_bank[3561],db_even.mem_bank[3561]);
$fdisplay(file, "0x1BD40,0x%h_0x%h", db_odd.mem_bank[3562],db_even.mem_bank[3562]);
$fdisplay(file, "0x1BD60,0x%h_0x%h", db_odd.mem_bank[3563],db_even.mem_bank[3563]);
$fdisplay(file, "0x1BD80,0x%h_0x%h", db_odd.mem_bank[3564],db_even.mem_bank[3564]);
$fdisplay(file, "0x1BDA0,0x%h_0x%h", db_odd.mem_bank[3565],db_even.mem_bank[3565]);
$fdisplay(file, "0x1BDC0,0x%h_0x%h", db_odd.mem_bank[3566],db_even.mem_bank[3566]);
$fdisplay(file, "0x1BDE0,0x%h_0x%h", db_odd.mem_bank[3567],db_even.mem_bank[3567]);
$fdisplay(file, "0x1BE00,0x%h_0x%h", db_odd.mem_bank[3568],db_even.mem_bank[3568]);
$fdisplay(file, "0x1BE20,0x%h_0x%h", db_odd.mem_bank[3569],db_even.mem_bank[3569]);
$fdisplay(file, "0x1BE40,0x%h_0x%h", db_odd.mem_bank[3570],db_even.mem_bank[3570]);
$fdisplay(file, "0x1BE60,0x%h_0x%h", db_odd.mem_bank[3571],db_even.mem_bank[3571]);
$fdisplay(file, "0x1BE80,0x%h_0x%h", db_odd.mem_bank[3572],db_even.mem_bank[3572]);
$fdisplay(file, "0x1BEA0,0x%h_0x%h", db_odd.mem_bank[3573],db_even.mem_bank[3573]);
$fdisplay(file, "0x1BEC0,0x%h_0x%h", db_odd.mem_bank[3574],db_even.mem_bank[3574]);
$fdisplay(file, "0x1BEE0,0x%h_0x%h", db_odd.mem_bank[3575],db_even.mem_bank[3575]);
$fdisplay(file, "0x1BF00,0x%h_0x%h", db_odd.mem_bank[3576],db_even.mem_bank[3576]);
$fdisplay(file, "0x1BF20,0x%h_0x%h", db_odd.mem_bank[3577],db_even.mem_bank[3577]);
$fdisplay(file, "0x1BF40,0x%h_0x%h", db_odd.mem_bank[3578],db_even.mem_bank[3578]);
$fdisplay(file, "0x1BF60,0x%h_0x%h", db_odd.mem_bank[3579],db_even.mem_bank[3579]);
$fdisplay(file, "0x1BF80,0x%h_0x%h", db_odd.mem_bank[3580],db_even.mem_bank[3580]);
$fdisplay(file, "0x1BFA0,0x%h_0x%h", db_odd.mem_bank[3581],db_even.mem_bank[3581]);
$fdisplay(file, "0x1BFC0,0x%h_0x%h", db_odd.mem_bank[3582],db_even.mem_bank[3582]);
$fdisplay(file, "0x1BFE0,0x%h_0x%h", db_odd.mem_bank[3583],db_even.mem_bank[3583]);
$fdisplay(file, "0x1C000,0x%h_0x%h", db_odd.mem_bank[3584],db_even.mem_bank[3584]);
$fdisplay(file, "0x1C020,0x%h_0x%h", db_odd.mem_bank[3585],db_even.mem_bank[3585]);
$fdisplay(file, "0x1C040,0x%h_0x%h", db_odd.mem_bank[3586],db_even.mem_bank[3586]);
$fdisplay(file, "0x1C060,0x%h_0x%h", db_odd.mem_bank[3587],db_even.mem_bank[3587]);
$fdisplay(file, "0x1C080,0x%h_0x%h", db_odd.mem_bank[3588],db_even.mem_bank[3588]);
$fdisplay(file, "0x1C0A0,0x%h_0x%h", db_odd.mem_bank[3589],db_even.mem_bank[3589]);
$fdisplay(file, "0x1C0C0,0x%h_0x%h", db_odd.mem_bank[3590],db_even.mem_bank[3590]);
$fdisplay(file, "0x1C0E0,0x%h_0x%h", db_odd.mem_bank[3591],db_even.mem_bank[3591]);
$fdisplay(file, "0x1C100,0x%h_0x%h", db_odd.mem_bank[3592],db_even.mem_bank[3592]);
$fdisplay(file, "0x1C120,0x%h_0x%h", db_odd.mem_bank[3593],db_even.mem_bank[3593]);
$fdisplay(file, "0x1C140,0x%h_0x%h", db_odd.mem_bank[3594],db_even.mem_bank[3594]);
$fdisplay(file, "0x1C160,0x%h_0x%h", db_odd.mem_bank[3595],db_even.mem_bank[3595]);
$fdisplay(file, "0x1C180,0x%h_0x%h", db_odd.mem_bank[3596],db_even.mem_bank[3596]);
$fdisplay(file, "0x1C1A0,0x%h_0x%h", db_odd.mem_bank[3597],db_even.mem_bank[3597]);
$fdisplay(file, "0x1C1C0,0x%h_0x%h", db_odd.mem_bank[3598],db_even.mem_bank[3598]);
$fdisplay(file, "0x1C1E0,0x%h_0x%h", db_odd.mem_bank[3599],db_even.mem_bank[3599]);
$fdisplay(file, "0x1C200,0x%h_0x%h", db_odd.mem_bank[3600],db_even.mem_bank[3600]);
$fdisplay(file, "0x1C220,0x%h_0x%h", db_odd.mem_bank[3601],db_even.mem_bank[3601]);
$fdisplay(file, "0x1C240,0x%h_0x%h", db_odd.mem_bank[3602],db_even.mem_bank[3602]);
$fdisplay(file, "0x1C260,0x%h_0x%h", db_odd.mem_bank[3603],db_even.mem_bank[3603]);
$fdisplay(file, "0x1C280,0x%h_0x%h", db_odd.mem_bank[3604],db_even.mem_bank[3604]);
$fdisplay(file, "0x1C2A0,0x%h_0x%h", db_odd.mem_bank[3605],db_even.mem_bank[3605]);
$fdisplay(file, "0x1C2C0,0x%h_0x%h", db_odd.mem_bank[3606],db_even.mem_bank[3606]);
$fdisplay(file, "0x1C2E0,0x%h_0x%h", db_odd.mem_bank[3607],db_even.mem_bank[3607]);
$fdisplay(file, "0x1C300,0x%h_0x%h", db_odd.mem_bank[3608],db_even.mem_bank[3608]);
$fdisplay(file, "0x1C320,0x%h_0x%h", db_odd.mem_bank[3609],db_even.mem_bank[3609]);
$fdisplay(file, "0x1C340,0x%h_0x%h", db_odd.mem_bank[3610],db_even.mem_bank[3610]);
$fdisplay(file, "0x1C360,0x%h_0x%h", db_odd.mem_bank[3611],db_even.mem_bank[3611]);
$fdisplay(file, "0x1C380,0x%h_0x%h", db_odd.mem_bank[3612],db_even.mem_bank[3612]);
$fdisplay(file, "0x1C3A0,0x%h_0x%h", db_odd.mem_bank[3613],db_even.mem_bank[3613]);
$fdisplay(file, "0x1C3C0,0x%h_0x%h", db_odd.mem_bank[3614],db_even.mem_bank[3614]);
$fdisplay(file, "0x1C3E0,0x%h_0x%h", db_odd.mem_bank[3615],db_even.mem_bank[3615]);
$fdisplay(file, "0x1C400,0x%h_0x%h", db_odd.mem_bank[3616],db_even.mem_bank[3616]);
$fdisplay(file, "0x1C420,0x%h_0x%h", db_odd.mem_bank[3617],db_even.mem_bank[3617]);
$fdisplay(file, "0x1C440,0x%h_0x%h", db_odd.mem_bank[3618],db_even.mem_bank[3618]);
$fdisplay(file, "0x1C460,0x%h_0x%h", db_odd.mem_bank[3619],db_even.mem_bank[3619]);
$fdisplay(file, "0x1C480,0x%h_0x%h", db_odd.mem_bank[3620],db_even.mem_bank[3620]);
$fdisplay(file, "0x1C4A0,0x%h_0x%h", db_odd.mem_bank[3621],db_even.mem_bank[3621]);
$fdisplay(file, "0x1C4C0,0x%h_0x%h", db_odd.mem_bank[3622],db_even.mem_bank[3622]);
$fdisplay(file, "0x1C4E0,0x%h_0x%h", db_odd.mem_bank[3623],db_even.mem_bank[3623]);
$fdisplay(file, "0x1C500,0x%h_0x%h", db_odd.mem_bank[3624],db_even.mem_bank[3624]);
$fdisplay(file, "0x1C520,0x%h_0x%h", db_odd.mem_bank[3625],db_even.mem_bank[3625]);
$fdisplay(file, "0x1C540,0x%h_0x%h", db_odd.mem_bank[3626],db_even.mem_bank[3626]);
$fdisplay(file, "0x1C560,0x%h_0x%h", db_odd.mem_bank[3627],db_even.mem_bank[3627]);
$fdisplay(file, "0x1C580,0x%h_0x%h", db_odd.mem_bank[3628],db_even.mem_bank[3628]);
$fdisplay(file, "0x1C5A0,0x%h_0x%h", db_odd.mem_bank[3629],db_even.mem_bank[3629]);
$fdisplay(file, "0x1C5C0,0x%h_0x%h", db_odd.mem_bank[3630],db_even.mem_bank[3630]);
$fdisplay(file, "0x1C5E0,0x%h_0x%h", db_odd.mem_bank[3631],db_even.mem_bank[3631]);
$fdisplay(file, "0x1C600,0x%h_0x%h", db_odd.mem_bank[3632],db_even.mem_bank[3632]);
$fdisplay(file, "0x1C620,0x%h_0x%h", db_odd.mem_bank[3633],db_even.mem_bank[3633]);
$fdisplay(file, "0x1C640,0x%h_0x%h", db_odd.mem_bank[3634],db_even.mem_bank[3634]);
$fdisplay(file, "0x1C660,0x%h_0x%h", db_odd.mem_bank[3635],db_even.mem_bank[3635]);
$fdisplay(file, "0x1C680,0x%h_0x%h", db_odd.mem_bank[3636],db_even.mem_bank[3636]);
$fdisplay(file, "0x1C6A0,0x%h_0x%h", db_odd.mem_bank[3637],db_even.mem_bank[3637]);
$fdisplay(file, "0x1C6C0,0x%h_0x%h", db_odd.mem_bank[3638],db_even.mem_bank[3638]);
$fdisplay(file, "0x1C6E0,0x%h_0x%h", db_odd.mem_bank[3639],db_even.mem_bank[3639]);
$fdisplay(file, "0x1C700,0x%h_0x%h", db_odd.mem_bank[3640],db_even.mem_bank[3640]);
$fdisplay(file, "0x1C720,0x%h_0x%h", db_odd.mem_bank[3641],db_even.mem_bank[3641]);
$fdisplay(file, "0x1C740,0x%h_0x%h", db_odd.mem_bank[3642],db_even.mem_bank[3642]);
$fdisplay(file, "0x1C760,0x%h_0x%h", db_odd.mem_bank[3643],db_even.mem_bank[3643]);
$fdisplay(file, "0x1C780,0x%h_0x%h", db_odd.mem_bank[3644],db_even.mem_bank[3644]);
$fdisplay(file, "0x1C7A0,0x%h_0x%h", db_odd.mem_bank[3645],db_even.mem_bank[3645]);
$fdisplay(file, "0x1C7C0,0x%h_0x%h", db_odd.mem_bank[3646],db_even.mem_bank[3646]);
$fdisplay(file, "0x1C7E0,0x%h_0x%h", db_odd.mem_bank[3647],db_even.mem_bank[3647]);
$fdisplay(file, "0x1C800,0x%h_0x%h", db_odd.mem_bank[3648],db_even.mem_bank[3648]);
$fdisplay(file, "0x1C820,0x%h_0x%h", db_odd.mem_bank[3649],db_even.mem_bank[3649]);
$fdisplay(file, "0x1C840,0x%h_0x%h", db_odd.mem_bank[3650],db_even.mem_bank[3650]);
$fdisplay(file, "0x1C860,0x%h_0x%h", db_odd.mem_bank[3651],db_even.mem_bank[3651]);
$fdisplay(file, "0x1C880,0x%h_0x%h", db_odd.mem_bank[3652],db_even.mem_bank[3652]);
$fdisplay(file, "0x1C8A0,0x%h_0x%h", db_odd.mem_bank[3653],db_even.mem_bank[3653]);
$fdisplay(file, "0x1C8C0,0x%h_0x%h", db_odd.mem_bank[3654],db_even.mem_bank[3654]);
$fdisplay(file, "0x1C8E0,0x%h_0x%h", db_odd.mem_bank[3655],db_even.mem_bank[3655]);
$fdisplay(file, "0x1C900,0x%h_0x%h", db_odd.mem_bank[3656],db_even.mem_bank[3656]);
$fdisplay(file, "0x1C920,0x%h_0x%h", db_odd.mem_bank[3657],db_even.mem_bank[3657]);
$fdisplay(file, "0x1C940,0x%h_0x%h", db_odd.mem_bank[3658],db_even.mem_bank[3658]);
$fdisplay(file, "0x1C960,0x%h_0x%h", db_odd.mem_bank[3659],db_even.mem_bank[3659]);
$fdisplay(file, "0x1C980,0x%h_0x%h", db_odd.mem_bank[3660],db_even.mem_bank[3660]);
$fdisplay(file, "0x1C9A0,0x%h_0x%h", db_odd.mem_bank[3661],db_even.mem_bank[3661]);
$fdisplay(file, "0x1C9C0,0x%h_0x%h", db_odd.mem_bank[3662],db_even.mem_bank[3662]);
$fdisplay(file, "0x1C9E0,0x%h_0x%h", db_odd.mem_bank[3663],db_even.mem_bank[3663]);
$fdisplay(file, "0x1CA00,0x%h_0x%h", db_odd.mem_bank[3664],db_even.mem_bank[3664]);
$fdisplay(file, "0x1CA20,0x%h_0x%h", db_odd.mem_bank[3665],db_even.mem_bank[3665]);
$fdisplay(file, "0x1CA40,0x%h_0x%h", db_odd.mem_bank[3666],db_even.mem_bank[3666]);
$fdisplay(file, "0x1CA60,0x%h_0x%h", db_odd.mem_bank[3667],db_even.mem_bank[3667]);
$fdisplay(file, "0x1CA80,0x%h_0x%h", db_odd.mem_bank[3668],db_even.mem_bank[3668]);
$fdisplay(file, "0x1CAA0,0x%h_0x%h", db_odd.mem_bank[3669],db_even.mem_bank[3669]);
$fdisplay(file, "0x1CAC0,0x%h_0x%h", db_odd.mem_bank[3670],db_even.mem_bank[3670]);
$fdisplay(file, "0x1CAE0,0x%h_0x%h", db_odd.mem_bank[3671],db_even.mem_bank[3671]);
$fdisplay(file, "0x1CB00,0x%h_0x%h", db_odd.mem_bank[3672],db_even.mem_bank[3672]);
$fdisplay(file, "0x1CB20,0x%h_0x%h", db_odd.mem_bank[3673],db_even.mem_bank[3673]);
$fdisplay(file, "0x1CB40,0x%h_0x%h", db_odd.mem_bank[3674],db_even.mem_bank[3674]);
$fdisplay(file, "0x1CB60,0x%h_0x%h", db_odd.mem_bank[3675],db_even.mem_bank[3675]);
$fdisplay(file, "0x1CB80,0x%h_0x%h", db_odd.mem_bank[3676],db_even.mem_bank[3676]);
$fdisplay(file, "0x1CBA0,0x%h_0x%h", db_odd.mem_bank[3677],db_even.mem_bank[3677]);
$fdisplay(file, "0x1CBC0,0x%h_0x%h", db_odd.mem_bank[3678],db_even.mem_bank[3678]);
$fdisplay(file, "0x1CBE0,0x%h_0x%h", db_odd.mem_bank[3679],db_even.mem_bank[3679]);
$fdisplay(file, "0x1CC00,0x%h_0x%h", db_odd.mem_bank[3680],db_even.mem_bank[3680]);
$fdisplay(file, "0x1CC20,0x%h_0x%h", db_odd.mem_bank[3681],db_even.mem_bank[3681]);
$fdisplay(file, "0x1CC40,0x%h_0x%h", db_odd.mem_bank[3682],db_even.mem_bank[3682]);
$fdisplay(file, "0x1CC60,0x%h_0x%h", db_odd.mem_bank[3683],db_even.mem_bank[3683]);
$fdisplay(file, "0x1CC80,0x%h_0x%h", db_odd.mem_bank[3684],db_even.mem_bank[3684]);
$fdisplay(file, "0x1CCA0,0x%h_0x%h", db_odd.mem_bank[3685],db_even.mem_bank[3685]);
$fdisplay(file, "0x1CCC0,0x%h_0x%h", db_odd.mem_bank[3686],db_even.mem_bank[3686]);
$fdisplay(file, "0x1CCE0,0x%h_0x%h", db_odd.mem_bank[3687],db_even.mem_bank[3687]);
$fdisplay(file, "0x1CD00,0x%h_0x%h", db_odd.mem_bank[3688],db_even.mem_bank[3688]);
$fdisplay(file, "0x1CD20,0x%h_0x%h", db_odd.mem_bank[3689],db_even.mem_bank[3689]);
$fdisplay(file, "0x1CD40,0x%h_0x%h", db_odd.mem_bank[3690],db_even.mem_bank[3690]);
$fdisplay(file, "0x1CD60,0x%h_0x%h", db_odd.mem_bank[3691],db_even.mem_bank[3691]);
$fdisplay(file, "0x1CD80,0x%h_0x%h", db_odd.mem_bank[3692],db_even.mem_bank[3692]);
$fdisplay(file, "0x1CDA0,0x%h_0x%h", db_odd.mem_bank[3693],db_even.mem_bank[3693]);
$fdisplay(file, "0x1CDC0,0x%h_0x%h", db_odd.mem_bank[3694],db_even.mem_bank[3694]);
$fdisplay(file, "0x1CDE0,0x%h_0x%h", db_odd.mem_bank[3695],db_even.mem_bank[3695]);
$fdisplay(file, "0x1CE00,0x%h_0x%h", db_odd.mem_bank[3696],db_even.mem_bank[3696]);
$fdisplay(file, "0x1CE20,0x%h_0x%h", db_odd.mem_bank[3697],db_even.mem_bank[3697]);
$fdisplay(file, "0x1CE40,0x%h_0x%h", db_odd.mem_bank[3698],db_even.mem_bank[3698]);
$fdisplay(file, "0x1CE60,0x%h_0x%h", db_odd.mem_bank[3699],db_even.mem_bank[3699]);
$fdisplay(file, "0x1CE80,0x%h_0x%h", db_odd.mem_bank[3700],db_even.mem_bank[3700]);
$fdisplay(file, "0x1CEA0,0x%h_0x%h", db_odd.mem_bank[3701],db_even.mem_bank[3701]);
$fdisplay(file, "0x1CEC0,0x%h_0x%h", db_odd.mem_bank[3702],db_even.mem_bank[3702]);
$fdisplay(file, "0x1CEE0,0x%h_0x%h", db_odd.mem_bank[3703],db_even.mem_bank[3703]);
$fdisplay(file, "0x1CF00,0x%h_0x%h", db_odd.mem_bank[3704],db_even.mem_bank[3704]);
$fdisplay(file, "0x1CF20,0x%h_0x%h", db_odd.mem_bank[3705],db_even.mem_bank[3705]);
$fdisplay(file, "0x1CF40,0x%h_0x%h", db_odd.mem_bank[3706],db_even.mem_bank[3706]);
$fdisplay(file, "0x1CF60,0x%h_0x%h", db_odd.mem_bank[3707],db_even.mem_bank[3707]);
$fdisplay(file, "0x1CF80,0x%h_0x%h", db_odd.mem_bank[3708],db_even.mem_bank[3708]);
$fdisplay(file, "0x1CFA0,0x%h_0x%h", db_odd.mem_bank[3709],db_even.mem_bank[3709]);
$fdisplay(file, "0x1CFC0,0x%h_0x%h", db_odd.mem_bank[3710],db_even.mem_bank[3710]);
$fdisplay(file, "0x1CFE0,0x%h_0x%h", db_odd.mem_bank[3711],db_even.mem_bank[3711]);
$fdisplay(file, "0x1D000,0x%h_0x%h", db_odd.mem_bank[3712],db_even.mem_bank[3712]);
$fdisplay(file, "0x1D020,0x%h_0x%h", db_odd.mem_bank[3713],db_even.mem_bank[3713]);
$fdisplay(file, "0x1D040,0x%h_0x%h", db_odd.mem_bank[3714],db_even.mem_bank[3714]);
$fdisplay(file, "0x1D060,0x%h_0x%h", db_odd.mem_bank[3715],db_even.mem_bank[3715]);
$fdisplay(file, "0x1D080,0x%h_0x%h", db_odd.mem_bank[3716],db_even.mem_bank[3716]);
$fdisplay(file, "0x1D0A0,0x%h_0x%h", db_odd.mem_bank[3717],db_even.mem_bank[3717]);
$fdisplay(file, "0x1D0C0,0x%h_0x%h", db_odd.mem_bank[3718],db_even.mem_bank[3718]);
$fdisplay(file, "0x1D0E0,0x%h_0x%h", db_odd.mem_bank[3719],db_even.mem_bank[3719]);
$fdisplay(file, "0x1D100,0x%h_0x%h", db_odd.mem_bank[3720],db_even.mem_bank[3720]);
$fdisplay(file, "0x1D120,0x%h_0x%h", db_odd.mem_bank[3721],db_even.mem_bank[3721]);
$fdisplay(file, "0x1D140,0x%h_0x%h", db_odd.mem_bank[3722],db_even.mem_bank[3722]);
$fdisplay(file, "0x1D160,0x%h_0x%h", db_odd.mem_bank[3723],db_even.mem_bank[3723]);
$fdisplay(file, "0x1D180,0x%h_0x%h", db_odd.mem_bank[3724],db_even.mem_bank[3724]);
$fdisplay(file, "0x1D1A0,0x%h_0x%h", db_odd.mem_bank[3725],db_even.mem_bank[3725]);
$fdisplay(file, "0x1D1C0,0x%h_0x%h", db_odd.mem_bank[3726],db_even.mem_bank[3726]);
$fdisplay(file, "0x1D1E0,0x%h_0x%h", db_odd.mem_bank[3727],db_even.mem_bank[3727]);
$fdisplay(file, "0x1D200,0x%h_0x%h", db_odd.mem_bank[3728],db_even.mem_bank[3728]);
$fdisplay(file, "0x1D220,0x%h_0x%h", db_odd.mem_bank[3729],db_even.mem_bank[3729]);
$fdisplay(file, "0x1D240,0x%h_0x%h", db_odd.mem_bank[3730],db_even.mem_bank[3730]);
$fdisplay(file, "0x1D260,0x%h_0x%h", db_odd.mem_bank[3731],db_even.mem_bank[3731]);
$fdisplay(file, "0x1D280,0x%h_0x%h", db_odd.mem_bank[3732],db_even.mem_bank[3732]);
$fdisplay(file, "0x1D2A0,0x%h_0x%h", db_odd.mem_bank[3733],db_even.mem_bank[3733]);
$fdisplay(file, "0x1D2C0,0x%h_0x%h", db_odd.mem_bank[3734],db_even.mem_bank[3734]);
$fdisplay(file, "0x1D2E0,0x%h_0x%h", db_odd.mem_bank[3735],db_even.mem_bank[3735]);
$fdisplay(file, "0x1D300,0x%h_0x%h", db_odd.mem_bank[3736],db_even.mem_bank[3736]);
$fdisplay(file, "0x1D320,0x%h_0x%h", db_odd.mem_bank[3737],db_even.mem_bank[3737]);
$fdisplay(file, "0x1D340,0x%h_0x%h", db_odd.mem_bank[3738],db_even.mem_bank[3738]);
$fdisplay(file, "0x1D360,0x%h_0x%h", db_odd.mem_bank[3739],db_even.mem_bank[3739]);
$fdisplay(file, "0x1D380,0x%h_0x%h", db_odd.mem_bank[3740],db_even.mem_bank[3740]);
$fdisplay(file, "0x1D3A0,0x%h_0x%h", db_odd.mem_bank[3741],db_even.mem_bank[3741]);
$fdisplay(file, "0x1D3C0,0x%h_0x%h", db_odd.mem_bank[3742],db_even.mem_bank[3742]);
$fdisplay(file, "0x1D3E0,0x%h_0x%h", db_odd.mem_bank[3743],db_even.mem_bank[3743]);
$fdisplay(file, "0x1D400,0x%h_0x%h", db_odd.mem_bank[3744],db_even.mem_bank[3744]);
$fdisplay(file, "0x1D420,0x%h_0x%h", db_odd.mem_bank[3745],db_even.mem_bank[3745]);
$fdisplay(file, "0x1D440,0x%h_0x%h", db_odd.mem_bank[3746],db_even.mem_bank[3746]);
$fdisplay(file, "0x1D460,0x%h_0x%h", db_odd.mem_bank[3747],db_even.mem_bank[3747]);
$fdisplay(file, "0x1D480,0x%h_0x%h", db_odd.mem_bank[3748],db_even.mem_bank[3748]);
$fdisplay(file, "0x1D4A0,0x%h_0x%h", db_odd.mem_bank[3749],db_even.mem_bank[3749]);
$fdisplay(file, "0x1D4C0,0x%h_0x%h", db_odd.mem_bank[3750],db_even.mem_bank[3750]);
$fdisplay(file, "0x1D4E0,0x%h_0x%h", db_odd.mem_bank[3751],db_even.mem_bank[3751]);
$fdisplay(file, "0x1D500,0x%h_0x%h", db_odd.mem_bank[3752],db_even.mem_bank[3752]);
$fdisplay(file, "0x1D520,0x%h_0x%h", db_odd.mem_bank[3753],db_even.mem_bank[3753]);
$fdisplay(file, "0x1D540,0x%h_0x%h", db_odd.mem_bank[3754],db_even.mem_bank[3754]);
$fdisplay(file, "0x1D560,0x%h_0x%h", db_odd.mem_bank[3755],db_even.mem_bank[3755]);
$fdisplay(file, "0x1D580,0x%h_0x%h", db_odd.mem_bank[3756],db_even.mem_bank[3756]);
$fdisplay(file, "0x1D5A0,0x%h_0x%h", db_odd.mem_bank[3757],db_even.mem_bank[3757]);
$fdisplay(file, "0x1D5C0,0x%h_0x%h", db_odd.mem_bank[3758],db_even.mem_bank[3758]);
$fdisplay(file, "0x1D5E0,0x%h_0x%h", db_odd.mem_bank[3759],db_even.mem_bank[3759]);
$fdisplay(file, "0x1D600,0x%h_0x%h", db_odd.mem_bank[3760],db_even.mem_bank[3760]);
$fdisplay(file, "0x1D620,0x%h_0x%h", db_odd.mem_bank[3761],db_even.mem_bank[3761]);
$fdisplay(file, "0x1D640,0x%h_0x%h", db_odd.mem_bank[3762],db_even.mem_bank[3762]);
$fdisplay(file, "0x1D660,0x%h_0x%h", db_odd.mem_bank[3763],db_even.mem_bank[3763]);
$fdisplay(file, "0x1D680,0x%h_0x%h", db_odd.mem_bank[3764],db_even.mem_bank[3764]);
$fdisplay(file, "0x1D6A0,0x%h_0x%h", db_odd.mem_bank[3765],db_even.mem_bank[3765]);
$fdisplay(file, "0x1D6C0,0x%h_0x%h", db_odd.mem_bank[3766],db_even.mem_bank[3766]);
$fdisplay(file, "0x1D6E0,0x%h_0x%h", db_odd.mem_bank[3767],db_even.mem_bank[3767]);
$fdisplay(file, "0x1D700,0x%h_0x%h", db_odd.mem_bank[3768],db_even.mem_bank[3768]);
$fdisplay(file, "0x1D720,0x%h_0x%h", db_odd.mem_bank[3769],db_even.mem_bank[3769]);
$fdisplay(file, "0x1D740,0x%h_0x%h", db_odd.mem_bank[3770],db_even.mem_bank[3770]);
$fdisplay(file, "0x1D760,0x%h_0x%h", db_odd.mem_bank[3771],db_even.mem_bank[3771]);
$fdisplay(file, "0x1D780,0x%h_0x%h", db_odd.mem_bank[3772],db_even.mem_bank[3772]);
$fdisplay(file, "0x1D7A0,0x%h_0x%h", db_odd.mem_bank[3773],db_even.mem_bank[3773]);
$fdisplay(file, "0x1D7C0,0x%h_0x%h", db_odd.mem_bank[3774],db_even.mem_bank[3774]);
$fdisplay(file, "0x1D7E0,0x%h_0x%h", db_odd.mem_bank[3775],db_even.mem_bank[3775]);
$fdisplay(file, "0x1D800,0x%h_0x%h", db_odd.mem_bank[3776],db_even.mem_bank[3776]);
$fdisplay(file, "0x1D820,0x%h_0x%h", db_odd.mem_bank[3777],db_even.mem_bank[3777]);
$fdisplay(file, "0x1D840,0x%h_0x%h", db_odd.mem_bank[3778],db_even.mem_bank[3778]);
$fdisplay(file, "0x1D860,0x%h_0x%h", db_odd.mem_bank[3779],db_even.mem_bank[3779]);
$fdisplay(file, "0x1D880,0x%h_0x%h", db_odd.mem_bank[3780],db_even.mem_bank[3780]);
$fdisplay(file, "0x1D8A0,0x%h_0x%h", db_odd.mem_bank[3781],db_even.mem_bank[3781]);
$fdisplay(file, "0x1D8C0,0x%h_0x%h", db_odd.mem_bank[3782],db_even.mem_bank[3782]);
$fdisplay(file, "0x1D8E0,0x%h_0x%h", db_odd.mem_bank[3783],db_even.mem_bank[3783]);
$fdisplay(file, "0x1D900,0x%h_0x%h", db_odd.mem_bank[3784],db_even.mem_bank[3784]);
$fdisplay(file, "0x1D920,0x%h_0x%h", db_odd.mem_bank[3785],db_even.mem_bank[3785]);
$fdisplay(file, "0x1D940,0x%h_0x%h", db_odd.mem_bank[3786],db_even.mem_bank[3786]);
$fdisplay(file, "0x1D960,0x%h_0x%h", db_odd.mem_bank[3787],db_even.mem_bank[3787]);
$fdisplay(file, "0x1D980,0x%h_0x%h", db_odd.mem_bank[3788],db_even.mem_bank[3788]);
$fdisplay(file, "0x1D9A0,0x%h_0x%h", db_odd.mem_bank[3789],db_even.mem_bank[3789]);
$fdisplay(file, "0x1D9C0,0x%h_0x%h", db_odd.mem_bank[3790],db_even.mem_bank[3790]);
$fdisplay(file, "0x1D9E0,0x%h_0x%h", db_odd.mem_bank[3791],db_even.mem_bank[3791]);
$fdisplay(file, "0x1DA00,0x%h_0x%h", db_odd.mem_bank[3792],db_even.mem_bank[3792]);
$fdisplay(file, "0x1DA20,0x%h_0x%h", db_odd.mem_bank[3793],db_even.mem_bank[3793]);
$fdisplay(file, "0x1DA40,0x%h_0x%h", db_odd.mem_bank[3794],db_even.mem_bank[3794]);
$fdisplay(file, "0x1DA60,0x%h_0x%h", db_odd.mem_bank[3795],db_even.mem_bank[3795]);
$fdisplay(file, "0x1DA80,0x%h_0x%h", db_odd.mem_bank[3796],db_even.mem_bank[3796]);
$fdisplay(file, "0x1DAA0,0x%h_0x%h", db_odd.mem_bank[3797],db_even.mem_bank[3797]);
$fdisplay(file, "0x1DAC0,0x%h_0x%h", db_odd.mem_bank[3798],db_even.mem_bank[3798]);
$fdisplay(file, "0x1DAE0,0x%h_0x%h", db_odd.mem_bank[3799],db_even.mem_bank[3799]);
$fdisplay(file, "0x1DB00,0x%h_0x%h", db_odd.mem_bank[3800],db_even.mem_bank[3800]);
$fdisplay(file, "0x1DB20,0x%h_0x%h", db_odd.mem_bank[3801],db_even.mem_bank[3801]);
$fdisplay(file, "0x1DB40,0x%h_0x%h", db_odd.mem_bank[3802],db_even.mem_bank[3802]);
$fdisplay(file, "0x1DB60,0x%h_0x%h", db_odd.mem_bank[3803],db_even.mem_bank[3803]);
$fdisplay(file, "0x1DB80,0x%h_0x%h", db_odd.mem_bank[3804],db_even.mem_bank[3804]);
$fdisplay(file, "0x1DBA0,0x%h_0x%h", db_odd.mem_bank[3805],db_even.mem_bank[3805]);
$fdisplay(file, "0x1DBC0,0x%h_0x%h", db_odd.mem_bank[3806],db_even.mem_bank[3806]);
$fdisplay(file, "0x1DBE0,0x%h_0x%h", db_odd.mem_bank[3807],db_even.mem_bank[3807]);
$fdisplay(file, "0x1DC00,0x%h_0x%h", db_odd.mem_bank[3808],db_even.mem_bank[3808]);
$fdisplay(file, "0x1DC20,0x%h_0x%h", db_odd.mem_bank[3809],db_even.mem_bank[3809]);
$fdisplay(file, "0x1DC40,0x%h_0x%h", db_odd.mem_bank[3810],db_even.mem_bank[3810]);
$fdisplay(file, "0x1DC60,0x%h_0x%h", db_odd.mem_bank[3811],db_even.mem_bank[3811]);
$fdisplay(file, "0x1DC80,0x%h_0x%h", db_odd.mem_bank[3812],db_even.mem_bank[3812]);
$fdisplay(file, "0x1DCA0,0x%h_0x%h", db_odd.mem_bank[3813],db_even.mem_bank[3813]);
$fdisplay(file, "0x1DCC0,0x%h_0x%h", db_odd.mem_bank[3814],db_even.mem_bank[3814]);
$fdisplay(file, "0x1DCE0,0x%h_0x%h", db_odd.mem_bank[3815],db_even.mem_bank[3815]);
$fdisplay(file, "0x1DD00,0x%h_0x%h", db_odd.mem_bank[3816],db_even.mem_bank[3816]);
$fdisplay(file, "0x1DD20,0x%h_0x%h", db_odd.mem_bank[3817],db_even.mem_bank[3817]);
$fdisplay(file, "0x1DD40,0x%h_0x%h", db_odd.mem_bank[3818],db_even.mem_bank[3818]);
$fdisplay(file, "0x1DD60,0x%h_0x%h", db_odd.mem_bank[3819],db_even.mem_bank[3819]);
$fdisplay(file, "0x1DD80,0x%h_0x%h", db_odd.mem_bank[3820],db_even.mem_bank[3820]);
$fdisplay(file, "0x1DDA0,0x%h_0x%h", db_odd.mem_bank[3821],db_even.mem_bank[3821]);
$fdisplay(file, "0x1DDC0,0x%h_0x%h", db_odd.mem_bank[3822],db_even.mem_bank[3822]);
$fdisplay(file, "0x1DDE0,0x%h_0x%h", db_odd.mem_bank[3823],db_even.mem_bank[3823]);
$fdisplay(file, "0x1DE00,0x%h_0x%h", db_odd.mem_bank[3824],db_even.mem_bank[3824]);
$fdisplay(file, "0x1DE20,0x%h_0x%h", db_odd.mem_bank[3825],db_even.mem_bank[3825]);
$fdisplay(file, "0x1DE40,0x%h_0x%h", db_odd.mem_bank[3826],db_even.mem_bank[3826]);
$fdisplay(file, "0x1DE60,0x%h_0x%h", db_odd.mem_bank[3827],db_even.mem_bank[3827]);
$fdisplay(file, "0x1DE80,0x%h_0x%h", db_odd.mem_bank[3828],db_even.mem_bank[3828]);
$fdisplay(file, "0x1DEA0,0x%h_0x%h", db_odd.mem_bank[3829],db_even.mem_bank[3829]);
$fdisplay(file, "0x1DEC0,0x%h_0x%h", db_odd.mem_bank[3830],db_even.mem_bank[3830]);
$fdisplay(file, "0x1DEE0,0x%h_0x%h", db_odd.mem_bank[3831],db_even.mem_bank[3831]);
$fdisplay(file, "0x1DF00,0x%h_0x%h", db_odd.mem_bank[3832],db_even.mem_bank[3832]);
$fdisplay(file, "0x1DF20,0x%h_0x%h", db_odd.mem_bank[3833],db_even.mem_bank[3833]);
$fdisplay(file, "0x1DF40,0x%h_0x%h", db_odd.mem_bank[3834],db_even.mem_bank[3834]);
$fdisplay(file, "0x1DF60,0x%h_0x%h", db_odd.mem_bank[3835],db_even.mem_bank[3835]);
$fdisplay(file, "0x1DF80,0x%h_0x%h", db_odd.mem_bank[3836],db_even.mem_bank[3836]);
$fdisplay(file, "0x1DFA0,0x%h_0x%h", db_odd.mem_bank[3837],db_even.mem_bank[3837]);
$fdisplay(file, "0x1DFC0,0x%h_0x%h", db_odd.mem_bank[3838],db_even.mem_bank[3838]);
$fdisplay(file, "0x1DFE0,0x%h_0x%h", db_odd.mem_bank[3839],db_even.mem_bank[3839]);
$fdisplay(file, "0x1E000,0x%h_0x%h", db_odd.mem_bank[3840],db_even.mem_bank[3840]);
$fdisplay(file, "0x1E020,0x%h_0x%h", db_odd.mem_bank[3841],db_even.mem_bank[3841]);
$fdisplay(file, "0x1E040,0x%h_0x%h", db_odd.mem_bank[3842],db_even.mem_bank[3842]);
$fdisplay(file, "0x1E060,0x%h_0x%h", db_odd.mem_bank[3843],db_even.mem_bank[3843]);
$fdisplay(file, "0x1E080,0x%h_0x%h", db_odd.mem_bank[3844],db_even.mem_bank[3844]);
$fdisplay(file, "0x1E0A0,0x%h_0x%h", db_odd.mem_bank[3845],db_even.mem_bank[3845]);
$fdisplay(file, "0x1E0C0,0x%h_0x%h", db_odd.mem_bank[3846],db_even.mem_bank[3846]);
$fdisplay(file, "0x1E0E0,0x%h_0x%h", db_odd.mem_bank[3847],db_even.mem_bank[3847]);
$fdisplay(file, "0x1E100,0x%h_0x%h", db_odd.mem_bank[3848],db_even.mem_bank[3848]);
$fdisplay(file, "0x1E120,0x%h_0x%h", db_odd.mem_bank[3849],db_even.mem_bank[3849]);
$fdisplay(file, "0x1E140,0x%h_0x%h", db_odd.mem_bank[3850],db_even.mem_bank[3850]);
$fdisplay(file, "0x1E160,0x%h_0x%h", db_odd.mem_bank[3851],db_even.mem_bank[3851]);
$fdisplay(file, "0x1E180,0x%h_0x%h", db_odd.mem_bank[3852],db_even.mem_bank[3852]);
$fdisplay(file, "0x1E1A0,0x%h_0x%h", db_odd.mem_bank[3853],db_even.mem_bank[3853]);
$fdisplay(file, "0x1E1C0,0x%h_0x%h", db_odd.mem_bank[3854],db_even.mem_bank[3854]);
$fdisplay(file, "0x1E1E0,0x%h_0x%h", db_odd.mem_bank[3855],db_even.mem_bank[3855]);
$fdisplay(file, "0x1E200,0x%h_0x%h", db_odd.mem_bank[3856],db_even.mem_bank[3856]);
$fdisplay(file, "0x1E220,0x%h_0x%h", db_odd.mem_bank[3857],db_even.mem_bank[3857]);
$fdisplay(file, "0x1E240,0x%h_0x%h", db_odd.mem_bank[3858],db_even.mem_bank[3858]);
$fdisplay(file, "0x1E260,0x%h_0x%h", db_odd.mem_bank[3859],db_even.mem_bank[3859]);
$fdisplay(file, "0x1E280,0x%h_0x%h", db_odd.mem_bank[3860],db_even.mem_bank[3860]);
$fdisplay(file, "0x1E2A0,0x%h_0x%h", db_odd.mem_bank[3861],db_even.mem_bank[3861]);
$fdisplay(file, "0x1E2C0,0x%h_0x%h", db_odd.mem_bank[3862],db_even.mem_bank[3862]);
$fdisplay(file, "0x1E2E0,0x%h_0x%h", db_odd.mem_bank[3863],db_even.mem_bank[3863]);
$fdisplay(file, "0x1E300,0x%h_0x%h", db_odd.mem_bank[3864],db_even.mem_bank[3864]);
$fdisplay(file, "0x1E320,0x%h_0x%h", db_odd.mem_bank[3865],db_even.mem_bank[3865]);
$fdisplay(file, "0x1E340,0x%h_0x%h", db_odd.mem_bank[3866],db_even.mem_bank[3866]);
$fdisplay(file, "0x1E360,0x%h_0x%h", db_odd.mem_bank[3867],db_even.mem_bank[3867]);
$fdisplay(file, "0x1E380,0x%h_0x%h", db_odd.mem_bank[3868],db_even.mem_bank[3868]);
$fdisplay(file, "0x1E3A0,0x%h_0x%h", db_odd.mem_bank[3869],db_even.mem_bank[3869]);
$fdisplay(file, "0x1E3C0,0x%h_0x%h", db_odd.mem_bank[3870],db_even.mem_bank[3870]);
$fdisplay(file, "0x1E3E0,0x%h_0x%h", db_odd.mem_bank[3871],db_even.mem_bank[3871]);
$fdisplay(file, "0x1E400,0x%h_0x%h", db_odd.mem_bank[3872],db_even.mem_bank[3872]);
$fdisplay(file, "0x1E420,0x%h_0x%h", db_odd.mem_bank[3873],db_even.mem_bank[3873]);
$fdisplay(file, "0x1E440,0x%h_0x%h", db_odd.mem_bank[3874],db_even.mem_bank[3874]);
$fdisplay(file, "0x1E460,0x%h_0x%h", db_odd.mem_bank[3875],db_even.mem_bank[3875]);
$fdisplay(file, "0x1E480,0x%h_0x%h", db_odd.mem_bank[3876],db_even.mem_bank[3876]);
$fdisplay(file, "0x1E4A0,0x%h_0x%h", db_odd.mem_bank[3877],db_even.mem_bank[3877]);
$fdisplay(file, "0x1E4C0,0x%h_0x%h", db_odd.mem_bank[3878],db_even.mem_bank[3878]);
$fdisplay(file, "0x1E4E0,0x%h_0x%h", db_odd.mem_bank[3879],db_even.mem_bank[3879]);
$fdisplay(file, "0x1E500,0x%h_0x%h", db_odd.mem_bank[3880],db_even.mem_bank[3880]);
$fdisplay(file, "0x1E520,0x%h_0x%h", db_odd.mem_bank[3881],db_even.mem_bank[3881]);
$fdisplay(file, "0x1E540,0x%h_0x%h", db_odd.mem_bank[3882],db_even.mem_bank[3882]);
$fdisplay(file, "0x1E560,0x%h_0x%h", db_odd.mem_bank[3883],db_even.mem_bank[3883]);
$fdisplay(file, "0x1E580,0x%h_0x%h", db_odd.mem_bank[3884],db_even.mem_bank[3884]);
$fdisplay(file, "0x1E5A0,0x%h_0x%h", db_odd.mem_bank[3885],db_even.mem_bank[3885]);
$fdisplay(file, "0x1E5C0,0x%h_0x%h", db_odd.mem_bank[3886],db_even.mem_bank[3886]);
$fdisplay(file, "0x1E5E0,0x%h_0x%h", db_odd.mem_bank[3887],db_even.mem_bank[3887]);
$fdisplay(file, "0x1E600,0x%h_0x%h", db_odd.mem_bank[3888],db_even.mem_bank[3888]);
$fdisplay(file, "0x1E620,0x%h_0x%h", db_odd.mem_bank[3889],db_even.mem_bank[3889]);
$fdisplay(file, "0x1E640,0x%h_0x%h", db_odd.mem_bank[3890],db_even.mem_bank[3890]);
$fdisplay(file, "0x1E660,0x%h_0x%h", db_odd.mem_bank[3891],db_even.mem_bank[3891]);
$fdisplay(file, "0x1E680,0x%h_0x%h", db_odd.mem_bank[3892],db_even.mem_bank[3892]);
$fdisplay(file, "0x1E6A0,0x%h_0x%h", db_odd.mem_bank[3893],db_even.mem_bank[3893]);
$fdisplay(file, "0x1E6C0,0x%h_0x%h", db_odd.mem_bank[3894],db_even.mem_bank[3894]);
$fdisplay(file, "0x1E6E0,0x%h_0x%h", db_odd.mem_bank[3895],db_even.mem_bank[3895]);
$fdisplay(file, "0x1E700,0x%h_0x%h", db_odd.mem_bank[3896],db_even.mem_bank[3896]);
$fdisplay(file, "0x1E720,0x%h_0x%h", db_odd.mem_bank[3897],db_even.mem_bank[3897]);
$fdisplay(file, "0x1E740,0x%h_0x%h", db_odd.mem_bank[3898],db_even.mem_bank[3898]);
$fdisplay(file, "0x1E760,0x%h_0x%h", db_odd.mem_bank[3899],db_even.mem_bank[3899]);
$fdisplay(file, "0x1E780,0x%h_0x%h", db_odd.mem_bank[3900],db_even.mem_bank[3900]);
$fdisplay(file, "0x1E7A0,0x%h_0x%h", db_odd.mem_bank[3901],db_even.mem_bank[3901]);
$fdisplay(file, "0x1E7C0,0x%h_0x%h", db_odd.mem_bank[3902],db_even.mem_bank[3902]);
$fdisplay(file, "0x1E7E0,0x%h_0x%h", db_odd.mem_bank[3903],db_even.mem_bank[3903]);
$fdisplay(file, "0x1E800,0x%h_0x%h", db_odd.mem_bank[3904],db_even.mem_bank[3904]);
$fdisplay(file, "0x1E820,0x%h_0x%h", db_odd.mem_bank[3905],db_even.mem_bank[3905]);
$fdisplay(file, "0x1E840,0x%h_0x%h", db_odd.mem_bank[3906],db_even.mem_bank[3906]);
$fdisplay(file, "0x1E860,0x%h_0x%h", db_odd.mem_bank[3907],db_even.mem_bank[3907]);
$fdisplay(file, "0x1E880,0x%h_0x%h", db_odd.mem_bank[3908],db_even.mem_bank[3908]);
$fdisplay(file, "0x1E8A0,0x%h_0x%h", db_odd.mem_bank[3909],db_even.mem_bank[3909]);
$fdisplay(file, "0x1E8C0,0x%h_0x%h", db_odd.mem_bank[3910],db_even.mem_bank[3910]);
$fdisplay(file, "0x1E8E0,0x%h_0x%h", db_odd.mem_bank[3911],db_even.mem_bank[3911]);
$fdisplay(file, "0x1E900,0x%h_0x%h", db_odd.mem_bank[3912],db_even.mem_bank[3912]);
$fdisplay(file, "0x1E920,0x%h_0x%h", db_odd.mem_bank[3913],db_even.mem_bank[3913]);
$fdisplay(file, "0x1E940,0x%h_0x%h", db_odd.mem_bank[3914],db_even.mem_bank[3914]);
$fdisplay(file, "0x1E960,0x%h_0x%h", db_odd.mem_bank[3915],db_even.mem_bank[3915]);
$fdisplay(file, "0x1E980,0x%h_0x%h", db_odd.mem_bank[3916],db_even.mem_bank[3916]);
$fdisplay(file, "0x1E9A0,0x%h_0x%h", db_odd.mem_bank[3917],db_even.mem_bank[3917]);
$fdisplay(file, "0x1E9C0,0x%h_0x%h", db_odd.mem_bank[3918],db_even.mem_bank[3918]);
$fdisplay(file, "0x1E9E0,0x%h_0x%h", db_odd.mem_bank[3919],db_even.mem_bank[3919]);
$fdisplay(file, "0x1EA00,0x%h_0x%h", db_odd.mem_bank[3920],db_even.mem_bank[3920]);
$fdisplay(file, "0x1EA20,0x%h_0x%h", db_odd.mem_bank[3921],db_even.mem_bank[3921]);
$fdisplay(file, "0x1EA40,0x%h_0x%h", db_odd.mem_bank[3922],db_even.mem_bank[3922]);
$fdisplay(file, "0x1EA60,0x%h_0x%h", db_odd.mem_bank[3923],db_even.mem_bank[3923]);
$fdisplay(file, "0x1EA80,0x%h_0x%h", db_odd.mem_bank[3924],db_even.mem_bank[3924]);
$fdisplay(file, "0x1EAA0,0x%h_0x%h", db_odd.mem_bank[3925],db_even.mem_bank[3925]);
$fdisplay(file, "0x1EAC0,0x%h_0x%h", db_odd.mem_bank[3926],db_even.mem_bank[3926]);
$fdisplay(file, "0x1EAE0,0x%h_0x%h", db_odd.mem_bank[3927],db_even.mem_bank[3927]);
$fdisplay(file, "0x1EB00,0x%h_0x%h", db_odd.mem_bank[3928],db_even.mem_bank[3928]);
$fdisplay(file, "0x1EB20,0x%h_0x%h", db_odd.mem_bank[3929],db_even.mem_bank[3929]);
$fdisplay(file, "0x1EB40,0x%h_0x%h", db_odd.mem_bank[3930],db_even.mem_bank[3930]);
$fdisplay(file, "0x1EB60,0x%h_0x%h", db_odd.mem_bank[3931],db_even.mem_bank[3931]);
$fdisplay(file, "0x1EB80,0x%h_0x%h", db_odd.mem_bank[3932],db_even.mem_bank[3932]);
$fdisplay(file, "0x1EBA0,0x%h_0x%h", db_odd.mem_bank[3933],db_even.mem_bank[3933]);
$fdisplay(file, "0x1EBC0,0x%h_0x%h", db_odd.mem_bank[3934],db_even.mem_bank[3934]);
$fdisplay(file, "0x1EBE0,0x%h_0x%h", db_odd.mem_bank[3935],db_even.mem_bank[3935]);
$fdisplay(file, "0x1EC00,0x%h_0x%h", db_odd.mem_bank[3936],db_even.mem_bank[3936]);
$fdisplay(file, "0x1EC20,0x%h_0x%h", db_odd.mem_bank[3937],db_even.mem_bank[3937]);
$fdisplay(file, "0x1EC40,0x%h_0x%h", db_odd.mem_bank[3938],db_even.mem_bank[3938]);
$fdisplay(file, "0x1EC60,0x%h_0x%h", db_odd.mem_bank[3939],db_even.mem_bank[3939]);
$fdisplay(file, "0x1EC80,0x%h_0x%h", db_odd.mem_bank[3940],db_even.mem_bank[3940]);
$fdisplay(file, "0x1ECA0,0x%h_0x%h", db_odd.mem_bank[3941],db_even.mem_bank[3941]);
$fdisplay(file, "0x1ECC0,0x%h_0x%h", db_odd.mem_bank[3942],db_even.mem_bank[3942]);
$fdisplay(file, "0x1ECE0,0x%h_0x%h", db_odd.mem_bank[3943],db_even.mem_bank[3943]);
$fdisplay(file, "0x1ED00,0x%h_0x%h", db_odd.mem_bank[3944],db_even.mem_bank[3944]);
$fdisplay(file, "0x1ED20,0x%h_0x%h", db_odd.mem_bank[3945],db_even.mem_bank[3945]);
$fdisplay(file, "0x1ED40,0x%h_0x%h", db_odd.mem_bank[3946],db_even.mem_bank[3946]);
$fdisplay(file, "0x1ED60,0x%h_0x%h", db_odd.mem_bank[3947],db_even.mem_bank[3947]);
$fdisplay(file, "0x1ED80,0x%h_0x%h", db_odd.mem_bank[3948],db_even.mem_bank[3948]);
$fdisplay(file, "0x1EDA0,0x%h_0x%h", db_odd.mem_bank[3949],db_even.mem_bank[3949]);
$fdisplay(file, "0x1EDC0,0x%h_0x%h", db_odd.mem_bank[3950],db_even.mem_bank[3950]);
$fdisplay(file, "0x1EDE0,0x%h_0x%h", db_odd.mem_bank[3951],db_even.mem_bank[3951]);
$fdisplay(file, "0x1EE00,0x%h_0x%h", db_odd.mem_bank[3952],db_even.mem_bank[3952]);
$fdisplay(file, "0x1EE20,0x%h_0x%h", db_odd.mem_bank[3953],db_even.mem_bank[3953]);
$fdisplay(file, "0x1EE40,0x%h_0x%h", db_odd.mem_bank[3954],db_even.mem_bank[3954]);
$fdisplay(file, "0x1EE60,0x%h_0x%h", db_odd.mem_bank[3955],db_even.mem_bank[3955]);
$fdisplay(file, "0x1EE80,0x%h_0x%h", db_odd.mem_bank[3956],db_even.mem_bank[3956]);
$fdisplay(file, "0x1EEA0,0x%h_0x%h", db_odd.mem_bank[3957],db_even.mem_bank[3957]);
$fdisplay(file, "0x1EEC0,0x%h_0x%h", db_odd.mem_bank[3958],db_even.mem_bank[3958]);
$fdisplay(file, "0x1EEE0,0x%h_0x%h", db_odd.mem_bank[3959],db_even.mem_bank[3959]);
$fdisplay(file, "0x1EF00,0x%h_0x%h", db_odd.mem_bank[3960],db_even.mem_bank[3960]);
$fdisplay(file, "0x1EF20,0x%h_0x%h", db_odd.mem_bank[3961],db_even.mem_bank[3961]);
$fdisplay(file, "0x1EF40,0x%h_0x%h", db_odd.mem_bank[3962],db_even.mem_bank[3962]);
$fdisplay(file, "0x1EF60,0x%h_0x%h", db_odd.mem_bank[3963],db_even.mem_bank[3963]);
$fdisplay(file, "0x1EF80,0x%h_0x%h", db_odd.mem_bank[3964],db_even.mem_bank[3964]);
$fdisplay(file, "0x1EFA0,0x%h_0x%h", db_odd.mem_bank[3965],db_even.mem_bank[3965]);
$fdisplay(file, "0x1EFC0,0x%h_0x%h", db_odd.mem_bank[3966],db_even.mem_bank[3966]);
$fdisplay(file, "0x1EFE0,0x%h_0x%h", db_odd.mem_bank[3967],db_even.mem_bank[3967]);
$fdisplay(file, "0x1F000,0x%h_0x%h", db_odd.mem_bank[3968],db_even.mem_bank[3968]);
$fdisplay(file, "0x1F020,0x%h_0x%h", db_odd.mem_bank[3969],db_even.mem_bank[3969]);
$fdisplay(file, "0x1F040,0x%h_0x%h", db_odd.mem_bank[3970],db_even.mem_bank[3970]);
$fdisplay(file, "0x1F060,0x%h_0x%h", db_odd.mem_bank[3971],db_even.mem_bank[3971]);
$fdisplay(file, "0x1F080,0x%h_0x%h", db_odd.mem_bank[3972],db_even.mem_bank[3972]);
$fdisplay(file, "0x1F0A0,0x%h_0x%h", db_odd.mem_bank[3973],db_even.mem_bank[3973]);
$fdisplay(file, "0x1F0C0,0x%h_0x%h", db_odd.mem_bank[3974],db_even.mem_bank[3974]);
$fdisplay(file, "0x1F0E0,0x%h_0x%h", db_odd.mem_bank[3975],db_even.mem_bank[3975]);
$fdisplay(file, "0x1F100,0x%h_0x%h", db_odd.mem_bank[3976],db_even.mem_bank[3976]);
$fdisplay(file, "0x1F120,0x%h_0x%h", db_odd.mem_bank[3977],db_even.mem_bank[3977]);
$fdisplay(file, "0x1F140,0x%h_0x%h", db_odd.mem_bank[3978],db_even.mem_bank[3978]);
$fdisplay(file, "0x1F160,0x%h_0x%h", db_odd.mem_bank[3979],db_even.mem_bank[3979]);
$fdisplay(file, "0x1F180,0x%h_0x%h", db_odd.mem_bank[3980],db_even.mem_bank[3980]);
$fdisplay(file, "0x1F1A0,0x%h_0x%h", db_odd.mem_bank[3981],db_even.mem_bank[3981]);
$fdisplay(file, "0x1F1C0,0x%h_0x%h", db_odd.mem_bank[3982],db_even.mem_bank[3982]);
$fdisplay(file, "0x1F1E0,0x%h_0x%h", db_odd.mem_bank[3983],db_even.mem_bank[3983]);
$fdisplay(file, "0x1F200,0x%h_0x%h", db_odd.mem_bank[3984],db_even.mem_bank[3984]);
$fdisplay(file, "0x1F220,0x%h_0x%h", db_odd.mem_bank[3985],db_even.mem_bank[3985]);
$fdisplay(file, "0x1F240,0x%h_0x%h", db_odd.mem_bank[3986],db_even.mem_bank[3986]);
$fdisplay(file, "0x1F260,0x%h_0x%h", db_odd.mem_bank[3987],db_even.mem_bank[3987]);
$fdisplay(file, "0x1F280,0x%h_0x%h", db_odd.mem_bank[3988],db_even.mem_bank[3988]);
$fdisplay(file, "0x1F2A0,0x%h_0x%h", db_odd.mem_bank[3989],db_even.mem_bank[3989]);
$fdisplay(file, "0x1F2C0,0x%h_0x%h", db_odd.mem_bank[3990],db_even.mem_bank[3990]);
$fdisplay(file, "0x1F2E0,0x%h_0x%h", db_odd.mem_bank[3991],db_even.mem_bank[3991]);
$fdisplay(file, "0x1F300,0x%h_0x%h", db_odd.mem_bank[3992],db_even.mem_bank[3992]);
$fdisplay(file, "0x1F320,0x%h_0x%h", db_odd.mem_bank[3993],db_even.mem_bank[3993]);
$fdisplay(file, "0x1F340,0x%h_0x%h", db_odd.mem_bank[3994],db_even.mem_bank[3994]);
$fdisplay(file, "0x1F360,0x%h_0x%h", db_odd.mem_bank[3995],db_even.mem_bank[3995]);
$fdisplay(file, "0x1F380,0x%h_0x%h", db_odd.mem_bank[3996],db_even.mem_bank[3996]);
$fdisplay(file, "0x1F3A0,0x%h_0x%h", db_odd.mem_bank[3997],db_even.mem_bank[3997]);
$fdisplay(file, "0x1F3C0,0x%h_0x%h", db_odd.mem_bank[3998],db_even.mem_bank[3998]);
$fdisplay(file, "0x1F3E0,0x%h_0x%h", db_odd.mem_bank[3999],db_even.mem_bank[3999]);
$fdisplay(file, "0x1F400,0x%h_0x%h", db_odd.mem_bank[4000],db_even.mem_bank[4000]);
$fdisplay(file, "0x1F420,0x%h_0x%h", db_odd.mem_bank[4001],db_even.mem_bank[4001]);
$fdisplay(file, "0x1F440,0x%h_0x%h", db_odd.mem_bank[4002],db_even.mem_bank[4002]);
$fdisplay(file, "0x1F460,0x%h_0x%h", db_odd.mem_bank[4003],db_even.mem_bank[4003]);
$fdisplay(file, "0x1F480,0x%h_0x%h", db_odd.mem_bank[4004],db_even.mem_bank[4004]);
$fdisplay(file, "0x1F4A0,0x%h_0x%h", db_odd.mem_bank[4005],db_even.mem_bank[4005]);
$fdisplay(file, "0x1F4C0,0x%h_0x%h", db_odd.mem_bank[4006],db_even.mem_bank[4006]);
$fdisplay(file, "0x1F4E0,0x%h_0x%h", db_odd.mem_bank[4007],db_even.mem_bank[4007]);
$fdisplay(file, "0x1F500,0x%h_0x%h", db_odd.mem_bank[4008],db_even.mem_bank[4008]);
$fdisplay(file, "0x1F520,0x%h_0x%h", db_odd.mem_bank[4009],db_even.mem_bank[4009]);
$fdisplay(file, "0x1F540,0x%h_0x%h", db_odd.mem_bank[4010],db_even.mem_bank[4010]);
$fdisplay(file, "0x1F560,0x%h_0x%h", db_odd.mem_bank[4011],db_even.mem_bank[4011]);
$fdisplay(file, "0x1F580,0x%h_0x%h", db_odd.mem_bank[4012],db_even.mem_bank[4012]);
$fdisplay(file, "0x1F5A0,0x%h_0x%h", db_odd.mem_bank[4013],db_even.mem_bank[4013]);
$fdisplay(file, "0x1F5C0,0x%h_0x%h", db_odd.mem_bank[4014],db_even.mem_bank[4014]);
$fdisplay(file, "0x1F5E0,0x%h_0x%h", db_odd.mem_bank[4015],db_even.mem_bank[4015]);
$fdisplay(file, "0x1F600,0x%h_0x%h", db_odd.mem_bank[4016],db_even.mem_bank[4016]);
$fdisplay(file, "0x1F620,0x%h_0x%h", db_odd.mem_bank[4017],db_even.mem_bank[4017]);
$fdisplay(file, "0x1F640,0x%h_0x%h", db_odd.mem_bank[4018],db_even.mem_bank[4018]);
$fdisplay(file, "0x1F660,0x%h_0x%h", db_odd.mem_bank[4019],db_even.mem_bank[4019]);
$fdisplay(file, "0x1F680,0x%h_0x%h", db_odd.mem_bank[4020],db_even.mem_bank[4020]);
$fdisplay(file, "0x1F6A0,0x%h_0x%h", db_odd.mem_bank[4021],db_even.mem_bank[4021]);
$fdisplay(file, "0x1F6C0,0x%h_0x%h", db_odd.mem_bank[4022],db_even.mem_bank[4022]);
$fdisplay(file, "0x1F6E0,0x%h_0x%h", db_odd.mem_bank[4023],db_even.mem_bank[4023]);
$fdisplay(file, "0x1F700,0x%h_0x%h", db_odd.mem_bank[4024],db_even.mem_bank[4024]);
$fdisplay(file, "0x1F720,0x%h_0x%h", db_odd.mem_bank[4025],db_even.mem_bank[4025]);
$fdisplay(file, "0x1F740,0x%h_0x%h", db_odd.mem_bank[4026],db_even.mem_bank[4026]);
$fdisplay(file, "0x1F760,0x%h_0x%h", db_odd.mem_bank[4027],db_even.mem_bank[4027]);
$fdisplay(file, "0x1F780,0x%h_0x%h", db_odd.mem_bank[4028],db_even.mem_bank[4028]);
$fdisplay(file, "0x1F7A0,0x%h_0x%h", db_odd.mem_bank[4029],db_even.mem_bank[4029]);
$fdisplay(file, "0x1F7C0,0x%h_0x%h", db_odd.mem_bank[4030],db_even.mem_bank[4030]);
$fdisplay(file, "0x1F7E0,0x%h_0x%h", db_odd.mem_bank[4031],db_even.mem_bank[4031]);
$fdisplay(file, "0x1F800,0x%h_0x%h", db_odd.mem_bank[4032],db_even.mem_bank[4032]);
$fdisplay(file, "0x1F820,0x%h_0x%h", db_odd.mem_bank[4033],db_even.mem_bank[4033]);
$fdisplay(file, "0x1F840,0x%h_0x%h", db_odd.mem_bank[4034],db_even.mem_bank[4034]);
$fdisplay(file, "0x1F860,0x%h_0x%h", db_odd.mem_bank[4035],db_even.mem_bank[4035]);
$fdisplay(file, "0x1F880,0x%h_0x%h", db_odd.mem_bank[4036],db_even.mem_bank[4036]);
$fdisplay(file, "0x1F8A0,0x%h_0x%h", db_odd.mem_bank[4037],db_even.mem_bank[4037]);
$fdisplay(file, "0x1F8C0,0x%h_0x%h", db_odd.mem_bank[4038],db_even.mem_bank[4038]);
$fdisplay(file, "0x1F8E0,0x%h_0x%h", db_odd.mem_bank[4039],db_even.mem_bank[4039]);
$fdisplay(file, "0x1F900,0x%h_0x%h", db_odd.mem_bank[4040],db_even.mem_bank[4040]);
$fdisplay(file, "0x1F920,0x%h_0x%h", db_odd.mem_bank[4041],db_even.mem_bank[4041]);
$fdisplay(file, "0x1F940,0x%h_0x%h", db_odd.mem_bank[4042],db_even.mem_bank[4042]);
$fdisplay(file, "0x1F960,0x%h_0x%h", db_odd.mem_bank[4043],db_even.mem_bank[4043]);
$fdisplay(file, "0x1F980,0x%h_0x%h", db_odd.mem_bank[4044],db_even.mem_bank[4044]);
$fdisplay(file, "0x1F9A0,0x%h_0x%h", db_odd.mem_bank[4045],db_even.mem_bank[4045]);
$fdisplay(file, "0x1F9C0,0x%h_0x%h", db_odd.mem_bank[4046],db_even.mem_bank[4046]);
$fdisplay(file, "0x1F9E0,0x%h_0x%h", db_odd.mem_bank[4047],db_even.mem_bank[4047]);
$fdisplay(file, "0x1FA00,0x%h_0x%h", db_odd.mem_bank[4048],db_even.mem_bank[4048]);
$fdisplay(file, "0x1FA20,0x%h_0x%h", db_odd.mem_bank[4049],db_even.mem_bank[4049]);
$fdisplay(file, "0x1FA40,0x%h_0x%h", db_odd.mem_bank[4050],db_even.mem_bank[4050]);
$fdisplay(file, "0x1FA60,0x%h_0x%h", db_odd.mem_bank[4051],db_even.mem_bank[4051]);
$fdisplay(file, "0x1FA80,0x%h_0x%h", db_odd.mem_bank[4052],db_even.mem_bank[4052]);
$fdisplay(file, "0x1FAA0,0x%h_0x%h", db_odd.mem_bank[4053],db_even.mem_bank[4053]);
$fdisplay(file, "0x1FAC0,0x%h_0x%h", db_odd.mem_bank[4054],db_even.mem_bank[4054]);
$fdisplay(file, "0x1FAE0,0x%h_0x%h", db_odd.mem_bank[4055],db_even.mem_bank[4055]);
$fdisplay(file, "0x1FB00,0x%h_0x%h", db_odd.mem_bank[4056],db_even.mem_bank[4056]);
$fdisplay(file, "0x1FB20,0x%h_0x%h", db_odd.mem_bank[4057],db_even.mem_bank[4057]);
$fdisplay(file, "0x1FB40,0x%h_0x%h", db_odd.mem_bank[4058],db_even.mem_bank[4058]);
$fdisplay(file, "0x1FB60,0x%h_0x%h", db_odd.mem_bank[4059],db_even.mem_bank[4059]);
$fdisplay(file, "0x1FB80,0x%h_0x%h", db_odd.mem_bank[4060],db_even.mem_bank[4060]);
$fdisplay(file, "0x1FBA0,0x%h_0x%h", db_odd.mem_bank[4061],db_even.mem_bank[4061]);
$fdisplay(file, "0x1FBC0,0x%h_0x%h", db_odd.mem_bank[4062],db_even.mem_bank[4062]);
$fdisplay(file, "0x1FBE0,0x%h_0x%h", db_odd.mem_bank[4063],db_even.mem_bank[4063]);
$fdisplay(file, "0x1FC00,0x%h_0x%h", db_odd.mem_bank[4064],db_even.mem_bank[4064]);
$fdisplay(file, "0x1FC20,0x%h_0x%h", db_odd.mem_bank[4065],db_even.mem_bank[4065]);
$fdisplay(file, "0x1FC40,0x%h_0x%h", db_odd.mem_bank[4066],db_even.mem_bank[4066]);
$fdisplay(file, "0x1FC60,0x%h_0x%h", db_odd.mem_bank[4067],db_even.mem_bank[4067]);
$fdisplay(file, "0x1FC80,0x%h_0x%h", db_odd.mem_bank[4068],db_even.mem_bank[4068]);
$fdisplay(file, "0x1FCA0,0x%h_0x%h", db_odd.mem_bank[4069],db_even.mem_bank[4069]);
$fdisplay(file, "0x1FCC0,0x%h_0x%h", db_odd.mem_bank[4070],db_even.mem_bank[4070]);
$fdisplay(file, "0x1FCE0,0x%h_0x%h", db_odd.mem_bank[4071],db_even.mem_bank[4071]);
$fdisplay(file, "0x1FD00,0x%h_0x%h", db_odd.mem_bank[4072],db_even.mem_bank[4072]);
$fdisplay(file, "0x1FD20,0x%h_0x%h", db_odd.mem_bank[4073],db_even.mem_bank[4073]);
$fdisplay(file, "0x1FD40,0x%h_0x%h", db_odd.mem_bank[4074],db_even.mem_bank[4074]);
$fdisplay(file, "0x1FD60,0x%h_0x%h", db_odd.mem_bank[4075],db_even.mem_bank[4075]);
$fdisplay(file, "0x1FD80,0x%h_0x%h", db_odd.mem_bank[4076],db_even.mem_bank[4076]);
$fdisplay(file, "0x1FDA0,0x%h_0x%h", db_odd.mem_bank[4077],db_even.mem_bank[4077]);
$fdisplay(file, "0x1FDC0,0x%h_0x%h", db_odd.mem_bank[4078],db_even.mem_bank[4078]);
$fdisplay(file, "0x1FDE0,0x%h_0x%h", db_odd.mem_bank[4079],db_even.mem_bank[4079]);
$fdisplay(file, "0x1FE00,0x%h_0x%h", db_odd.mem_bank[4080],db_even.mem_bank[4080]);
$fdisplay(file, "0x1FE20,0x%h_0x%h", db_odd.mem_bank[4081],db_even.mem_bank[4081]);
$fdisplay(file, "0x1FE40,0x%h_0x%h", db_odd.mem_bank[4082],db_even.mem_bank[4082]);
$fdisplay(file, "0x1FE60,0x%h_0x%h", db_odd.mem_bank[4083],db_even.mem_bank[4083]);
$fdisplay(file, "0x1FE80,0x%h_0x%h", db_odd.mem_bank[4084],db_even.mem_bank[4084]);
$fdisplay(file, "0x1FEA0,0x%h_0x%h", db_odd.mem_bank[4085],db_even.mem_bank[4085]);
$fdisplay(file, "0x1FEC0,0x%h_0x%h", db_odd.mem_bank[4086],db_even.mem_bank[4086]);
$fdisplay(file, "0x1FEE0,0x%h_0x%h", db_odd.mem_bank[4087],db_even.mem_bank[4087]);
$fdisplay(file, "0x1FF00,0x%h_0x%h", db_odd.mem_bank[4088],db_even.mem_bank[4088]);
$fdisplay(file, "0x1FF20,0x%h_0x%h", db_odd.mem_bank[4089],db_even.mem_bank[4089]);
$fdisplay(file, "0x1FF40,0x%h_0x%h", db_odd.mem_bank[4090],db_even.mem_bank[4090]);
$fdisplay(file, "0x1FF60,0x%h_0x%h", db_odd.mem_bank[4091],db_even.mem_bank[4091]);
$fdisplay(file, "0x1FF80,0x%h_0x%h", db_odd.mem_bank[4092],db_even.mem_bank[4092]);
$fdisplay(file, "0x1FFA0,0x%h_0x%h", db_odd.mem_bank[4093],db_even.mem_bank[4093]);
$fdisplay(file, "0x1FFC0,0x%h_0x%h", db_odd.mem_bank[4094],db_even.mem_bank[4094]);
$fdisplay(file, "0x1FFE0,0x%h_0x%h", db_odd.mem_bank[4095],db_even.mem_bank[4095]);

  end


endmodule